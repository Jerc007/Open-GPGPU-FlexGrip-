library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_reci is
	generic(
		word_bits	:natural:=13;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_reci is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1111110100000",
		"1111011100000",
		"1111000110000",
		"1110110000000",
		"1110011011000",
		"1110000110000",
		"1101110010000",
		"1101011111000",
		"1101001100000",
		"1100111010000",
		"1100101000000",
		"1100010111000",
		"1100000110000",
		"1011110101000",
		"1011100110000",
		"1011010110000",
		"1011000111000",
		"1010111001000",
		"1010101011000",
		"1010011101000",
		"1010001111000",
		"1010000010000",
		"1001110101000",
		"1001101001000",
		"1001011101000",
		"1001010001000",
		"1001000110000",
		"1000111011000",
		"1000110000000",
		"1000100101000",
		"1000011011000",
		"1000010001000",
		"1000000111000",
		"0111111101000",
		"0111110100000",
		"0111101011000",
		"0111100010000",
		"0111011001000",
		"0111010001000",
		"0111001000000",
		"0111000000000",
		"0110111000000",
		"0110110001000",
		"0110101001000",
		"0110100010000",
		"0110011011000",
		"0110010100000",
		"0110001101000",
		"0110000110000",
		"0110000000000",
		"0101111001000",
		"0101110011000",
		"0101101101000",
		"0101100111000",
		"0101100001000",
		"0101011011000",
		"0101010101000",
		"0101010000000",
		"0101001011000",
		"0101000101000",
		"0101000000000",
		"0100111011000",
		"0100110110000",
		"0100110001000",
		"0100101101000",
		"0100101000000",
		"0100100011000",
		"0100011111000",
		"0100011011000",
		"0100010110000",
		"0100010010000",
		"0100001110000",
		"0100001010000",
		"0100000110000",
		"0100000010000",
		"0011111110000",
		"0011111011000",
		"0011110111000",
		"0011110011000",
		"0011110000000",
		"0011101100000",
		"0011101001000",
		"0011100110000",
		"0011100010000",
		"0011011111000",
		"0011011100000",
		"0011011001000",
		"0011010110000",
		"0011010011000",
		"0011010000000",
		"0011001101000",
		"0011001011000",
		"0011001000000",
		"0011000101000",
		"0011000010000",
		"0011000000000",
		"0010111101000",
		"0010111011000",
		"0010111000000",
		"0010110110000",
		"0010110100000",
		"0010110001000",
		"0010101111000",
		"0010101101000",
		"0010101010000",
		"0010101000000",
		"0010100110000",
		"0010100100000",
		"0010100010000",
		"0010100000000",
		"0010011110000",
		"0010011100000",
		"0010011010000",
		"0010011000000",
		"0010010110000",
		"0010010100000",
		"0010010010000",
		"0010010001000",
		"0010001111000",
		"0010001101000",
		"0010001011000",
		"0010001010000",
		"0010001000000",
		"0010000110000",
		"0010000101000",
		"0010000011000",
		"0010000010000",
		"0010000000000"
	);
begin
	data <= "0"&rom(to_integer(unsigned(addr)));
end architecture;