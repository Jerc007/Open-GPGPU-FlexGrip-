library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci is
	generic(
		word_bits	:natural:=18;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"111111111111110100",
		"111111000000100100",
		"111110000010110000",
		"111101000110011000",
		"111100001011011000",
		"111011010001101100",
		"111010011001010000",
		"111001100010001000",
		"111000101100001000",
		"110111110111011000",
		"110111000011110000",
		"110110010001010000",
		"110101011111110100",
		"110100101111011000",
		"110100000000000000",
		"110011010001101000",
		"110010100100010000",
		"110001110111110000",
		"110001001100001100",
		"110000100001100000",
		"101111110111101100",
		"101111001110101100",
		"101110100110100000",
		"101101111111001000",
		"101101011000100100",
		"101100110010101100",
		"101100001101100100",
		"101011101001001100",
		"101011000101100000",
		"101010100010100000",
		"101010000000001000",
		"101001011110011100",
		"101000111101011000",
		"101000011100111000",
		"100111111101000000",
		"100111011101110000",
		"100110111111000100",
		"100110100000111000",
		"100110000011010100",
		"100101100110001100",
		"100101001001101000",
		"100100101101100100",
		"100100010010000000",
		"100011110110111100",
		"100011011100010100",
		"100011000010001100",
		"100010101000100000",
		"100010001111010000",
		"100001110110011100",
		"100001011110000000",
		"100001000110000000",
		"100000101110011000",
		"100000010111001100",
		"100000000000011000",
		"011111101001111100",
		"011111010011110100",
		"011110111110001000",
		"011110101000110000",
		"011110010011110000",
		"011101111111000100",
		"011101101010101100",
		"011101010110101000",
		"011101000010111100",
		"011100101111100000",
		"011100011100011000",
		"011100001001100100",
		"011011110111000100",
		"011011100100110100",
		"011011010010110100",
		"011011000001001000",
		"011010101111110000",
		"011010011110100100",
		"011010001101101100",
		"011001111101000000",
		"011001101100101000",
		"011001011100011100",
		"011001001100100000",
		"011000111100110100",
		"011000101101011000",
		"011000011110001000",
		"011000001111001000",
		"011000000000010100",
		"010111110001101100",
		"010111100011010100",
		"010111010101001000",
		"010111000111001000",
		"010110111001010100",
		"010110101011110000",
		"010110011110010100",
		"010110010001001000",
		"010110000100000100",
		"010101110111001100",
		"010101101010100000",
		"010101011110000000",
		"010101010001101000",
		"010101000101011100",
		"010100111001011100",
		"010100101101100100",
		"010100100001111000",
		"010100010110010100",
		"010100001010111100",
		"010011111111101100",
		"010011110100100100",
		"010011101001101000",
		"010011011110110000",
		"010011010100001000",
		"010011001001100100",
		"010010111111001000",
		"010010110100111000",
		"010010101010110000",
		"010010100000101100",
		"010010010110110100",
		"010010001101000100",
		"010010000011011000",
		"010001111001111000",
		"010001110000011100",
		"010001100111001000",
		"010001011110000000",
		"010001010100111000",
		"010001001011111100",
		"010001000011000100",
		"010000111010010100",
		"010000110001101100",
		"010000101001001100",
		"010000100000110000",
		"010000011000011000",
		"010000010000001000",
		"010000001000000000"
	);
begin
	data <= "10"&rom(to_integer(unsigned(addr)));
end architecture;