library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_sqrt_2_4 is
	generic(
		word_bits	:natural:=27;
		bus_bits	:natural:=29;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"011010100000100111100110100",
		"011011001101101100101011100",
		"011011111010011011101010000",
		"011100100110110101000001100",
		"011101010010111001010001000",
		"011101111110101000110101100",
		"011110101010000100001101000",
		"011111010101001011110010000",
		"100000000000000000000000000",
		"100000101010100001010000000",
		"100001010100101111111011000",
		"100001111110101100011001100",
		"100010101000010111000010000",
		"100011010001110000001100000",
		"100011111010111000001100000",
		"100100100011101111010111100",
		"100101001100010110000011100",
		"100101110100101100100011000",
		"100110011100110011001001100",
		"100111000100101010001001000",
		"100111101100010001110100100",
		"101000010011101010011100100",
		"101000111010110100010010100",
		"101001100001101111100110100",
		"101010001000011100101001000",
		"101010101110111011101001100",
		"101011010101001100110110100",
		"101011111011010000011111000",
		"101100100001000110110001100",
		"101101000110101111111100000",
		"101101101100001100001011100",
		"101110010001011011101101000",
		"101110110110011110101110100",
		"101111011011010101011011000",
		"110000000000000000000000000",
		"110000100100011110101000000",
		"110001001000110001100000000",
		"110001101100111000110010000",
		"110010010000110100101001100",
		"110010110100100101010001100",
		"110011011000001010110100000",
		"110011111011100101011011100",
		"110100011110110101010010000",
		"110101000001111010100000100",
		"110101100100110101010001100",
		"110110000111100101101110000",
		"110110101010001011111111000",
		"110111001100101000001101000",
		"110111101110111010100001000",
		"111000010001000011000011100",
		"111000110011000001111100100",
		"111001010100110111010100100",
		"111001110110100011010011100",
		"111010011000000110000000100",
		"111010111001011111100100000",
		"111011011010110000000101000",
		"111011111011110111101011000",
		"111100011100110110011100100",
		"111100111101101100100001000",
		"111101011110011001111111100",
		"111101111110111110111110100",
		"111110011111011011100100100",
		"111110111111101111110111100",
		"111111011111111011111111000"
	);
begin
	data <= "01"&rom(to_integer(unsigned(addr)));
end architecture;