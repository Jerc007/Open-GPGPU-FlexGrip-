
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TP_instructions is
	port(
		instruction_pointer_in : in  integer;
		num_instructions_out   : out integer;
		instruction_out        : out std_logic_vector(31 downto 0)
	);
end TP_instructions;

architecture arch of TP_instructions is
	constant TP_INSTRUCTIONS : integer := 726;

begin
	num_instructions_out <= TP_INSTRUCTIONS;

	process(instruction_pointer_in)
	begin
		case instruction_pointer_in is
			when 0 => instruction_out <= x"a000440d";   -- I2I.U32.U16 R3, g [0x2].U16;
when 1 => instruction_out <= x"04200780";
when 2 => instruction_out <= x"a0004215";   -- I2I.U32.U16 R5, g [0x1].U16;
when 3 => instruction_out <= x"04200780";
when 4 => instruction_out <= x"400b0c05";   -- IMUL.U16.U16 R1, R3L, R5H;
when 5 => instruction_out <= x"00000780";
when 6 => instruction_out <= x"600a0e05";   -- IMAD.U16 R1, R3H, R5L, R1;
when 7 => instruction_out <= x"00004780";
when 8 => instruction_out <= x"30100205";   -- SHL R1, R1, 0x10;
when 9 => instruction_out <= x"c4100780";
when 10 => instruction_out <= x"a0004619";   -- I2I.U32.U16 R6, g [0x3].U16;
when 11 => instruction_out <= x"04200780";
when 12 => instruction_out <= x"600a0c05";   -- IMAD.U16 R1, R3L, R5L, R1;
when 13 => instruction_out <= x"00004780";
when 14 => instruction_out <= x"400d0409";   -- IMUL.U16.U16 R2, R1L, R6H;
when 15 => instruction_out <= x"00000780";
when 16 => instruction_out <= x"600c0609";   -- IMAD.U16 R2, R1H, R6L, R2;
when 17 => instruction_out <= x"00008780";
when 18 => instruction_out <= x"30100409";   -- SHL R2, R2, 0x10;
when 19 => instruction_out <= x"c4100780";
when 20 => instruction_out <= x"600c0405";   -- IMAD.U16 R1, R1L, R6L, R2;
when 21 => instruction_out <= x"00008780";
when 22 => instruction_out <= x"a0004811";   -- I2I.U32.U16 R4, g [0x4].U16;
when 23 => instruction_out <= x"04200780";
when 24 => instruction_out <= x"40090409";   -- IMUL.U16.U16 R2, R1L, R4H;
when 25 => instruction_out <= x"00000780";
when 26 => instruction_out <= x"60080609";   -- IMAD.U16 R2, R1H, R4L, R2;
when 27 => instruction_out <= x"00008780";
when 28 => instruction_out <= x"30100409";   -- SHL R2, R2, 0x10;
when 29 => instruction_out <= x"c4100780";
when 30 => instruction_out <= x"60080421";   -- IMAD.U16 R8, R1L, R4L, R2;
when 31 => instruction_out <= x"00008780";
when 32 => instruction_out <= x"1100ee04";   -- MOV32 R1, g [0x7];
when 33 => instruction_out <= x"1100ec08";   -- MOV32 R2, g [0x6];
when 34 => instruction_out <= x"a0004a1d";   -- I2I.U32.U16 R7, g [0x5].U16;
when 35 => instruction_out <= x"04200780";
when 36 => instruction_out <= x"40050424";   -- IMUL32.U16.U16 R9, R1L, R2H;
when 37 => instruction_out <= x"40111c28";   -- IMUL32.U16.U16 R10, R7L, R8H;
when 38 => instruction_out <= x"60040625";   -- IMAD.U16 R9, R1H, R2L, R9;
when 39 => instruction_out <= x"00024780";
when 40 => instruction_out <= x"60101e29";   -- IMAD.U16 R10, R7H, R8L, R10;
when 41 => instruction_out <= x"00028780";
when 42 => instruction_out <= x"30101225";   -- SHL R9, R9, 0x10;
when 43 => instruction_out <= x"c4100780";
when 44 => instruction_out <= x"30101429";   -- SHL R10, R10, 0x10;
when 45 => instruction_out <= x"c4100780";
when 46 => instruction_out <= x"60040409";   -- IMAD.U16 R2, R1L, R2L, R9;
when 47 => instruction_out <= x"00024780";
when 48 => instruction_out <= x"60101c05";   -- IMAD.U16 R1, R7L, R8L, R10;
when 49 => instruction_out <= x"00028780";
when 50 => instruction_out <= x"307c05fd";   -- ISET.S32.C0 o[0x7f], R2, R124, LE;
when 51 => instruction_out <= x"6c00c7c8";
when 52 => instruction_out <= x"10021003";   -- BRA C0.NE, 0x108;
when 53 => instruction_out <= x"00000280";
when 54 => instruction_out <= x"1000f821";   -- MOV R8, R124;
when 55 => instruction_out <= x"0403c780";
when 56 => instruction_out <= x"30010409";   -- SHR.S32 R2, R2, 0x1;
when 57 => instruction_out <= x"ec100780";
when 58 => instruction_out <= x"307c05fd";   -- ISET.S32.C0 o[0x7f], R2, R124, GT;
when 59 => instruction_out <= x"6c0107c8";
when 60 => instruction_out <= x"20019021";   -- IADD32I R8, R8, 0x1;
when 61 => instruction_out <= x"00000003";
when 62 => instruction_out <= x"1001c003";   -- BRA C0.NE, 0xe0;
when 63 => instruction_out <= x"00000280";
when 64 => instruction_out <= x"10022003";   -- BRA  0x110;
when 65 => instruction_out <= x"00000780";
when 66 => instruction_out <= x"1000f821";   -- MOV R8, R124;
when 67 => instruction_out <= x"0403c780";
when 68 => instruction_out <= x"307c03fd";   -- ISET.S32.C0 o[0x7f], R1, R124, LE;
when 69 => instruction_out <= x"6c00c7c8";
when 70 => instruction_out <= x"1002a003";   -- BRA C0.NE, 0x150;
when 71 => instruction_out <= x"00000280";
when 72 => instruction_out <= x"1000f825";   -- MOV R9, R124;
when 73 => instruction_out <= x"0403c780";
when 74 => instruction_out <= x"30010205";   -- SHR.S32 R1, R1, 0x1;
when 75 => instruction_out <= x"ec100780";
when 76 => instruction_out <= x"307c03fd";   -- ISET.S32.C0 o[0x7f], R1, R124, GT;
when 77 => instruction_out <= x"6c0107c8";
when 78 => instruction_out <= x"20019225";   -- IADD32I R9, R9, 0x1;
when 79 => instruction_out <= x"00000003";
when 80 => instruction_out <= x"10025003";   -- BRA C0.NE, 0x128;
when 81 => instruction_out <= x"00000280";
when 82 => instruction_out <= x"1002b003";   -- BRA  0x158;
when 83 => instruction_out <= x"00000780";
when 84 => instruction_out <= x"1000f825";   -- MOV R9, R124;
when 85 => instruction_out <= x"0403c780";
when 86 => instruction_out <= x"a0004e05";   -- I2I.U32.U16 R1, g [0x7].U16;
when 87 => instruction_out <= x"04200780";
when 88 => instruction_out <= x"40021609";   -- IMUL.U16.U16 R2, R5H, R1L;
when 89 => instruction_out <= x"00000780";
when 90 => instruction_out <= x"60031409";   -- IMAD.U16 R2, R5L, R1H, R2;
when 91 => instruction_out <= x"00008780";
when 92 => instruction_out <= x"30100409";   -- SHL R2, R2, 0x10;
when 93 => instruction_out <= x"c4100780";
when 94 => instruction_out <= x"60021405";   -- IMAD.U16 R1, R5L, R1L, R2;
when 95 => instruction_out <= x"00008780";
when 96 => instruction_out <= x"a0004c1d";   -- I2I.U32.U16 R7, g [0x6].U16;
when 97 => instruction_out <= x"04200780";
when 98 => instruction_out <= x"300a0211";   -- SHR.U16 R2L, R0H, 0xa;
when 99 => instruction_out <= x"e0100780";
when 100 => instruction_out <= x"400e1628";   -- IMUL32.U16.U16 R10, R5H, R7L;
when 101 => instruction_out <= x"40020e2c";   -- IMUL32.U16.U16 R11, R3H, R1L;
when 102 => instruction_out <= x"a0000809";   -- I2I.U32.U16 R2, R2L;
when 103 => instruction_out <= x"04000780";
when 104 => instruction_out <= x"600f1429";   -- IMAD.U16 R10, R5L, R7H, R10;
when 105 => instruction_out <= x"00028780";
when 106 => instruction_out <= x"60030c31";   -- IMAD.U16 R12, R3L, R1H, R11;
when 107 => instruction_out <= x"0002c780";
when 108 => instruction_out <= x"20499024";   -- IADD32 R9, R8, -R9;
when 109 => instruction_out <= x"40041620";   -- IMUL32.U16.U16 R8, R5H, R2L;
when 110 => instruction_out <= x"3010142d";   -- SHL R11, R10, 0x10;
when 111 => instruction_out <= x"c4100780";
when 112 => instruction_out <= x"30101831";   -- SHL R12, R12, 0x10;
when 113 => instruction_out <= x"c4100780";
when 114 => instruction_out <= x"d0800205";   -- LOP.AND.U16 R0H, R0H, c[0x1][0x0];
when 115 => instruction_out <= x"00400780";
when 116 => instruction_out <= x"60051429";   -- IMAD.U16 R10, R5L, R2H, R8;
when 117 => instruction_out <= x"00020780";
when 118 => instruction_out <= x"600e141d";   -- IMAD.U16 R7, R5L, R7L, R11;
when 119 => instruction_out <= x"0002c780";
when 120 => instruction_out <= x"60020c21";   -- IMAD.U16 R8, R3L, R1L, R12;
when 121 => instruction_out <= x"00030780";
when 122 => instruction_out <= x"a0000205";   -- I2I.U32.U16 R1, R0H;
when 123 => instruction_out <= x"04000780";
when 124 => instruction_out <= x"3010142d";   -- SHL R11, R10, 0x10;
when 125 => instruction_out <= x"c4100780";
when 126 => instruction_out <= x"400b0429";   -- IMUL.U16.U16 R10, R1L, R5H;
when 127 => instruction_out <= x"00000780";
when 128 => instruction_out <= x"60041409";   -- IMAD.U16 R2, R5L, R2L, R11;
when 129 => instruction_out <= x"0002c780";
when 130 => instruction_out <= x"400e0e2d";   -- IMUL.U16.U16 R11, R3H, R7L;
when 131 => instruction_out <= x"00000780";
when 132 => instruction_out <= x"600a0629";   -- IMAD.U16 R10, R1H, R5L, R10;
when 133 => instruction_out <= x"00028780";
when 134 => instruction_out <= x"40101a35";   -- IMUL.U16.U16 R13, R6H, R8L;
when 135 => instruction_out <= x"00000780";
when 136 => instruction_out <= x"600f0c31";   -- IMAD.U16 R12, R3L, R7H, R11;
when 137 => instruction_out <= x"0002c780";
when 138 => instruction_out <= x"30101429";   -- SHL R10, R10, 0x10;
when 139 => instruction_out <= x"c4100780";
when 140 => instruction_out <= x"60111835";   -- IMAD.U16 R13, R6L, R8H, R13;
when 141 => instruction_out <= x"00034780";
when 142 => instruction_out <= x"4007082d";   -- IMUL.U16.U16 R11, R2L, R3H;
when 143 => instruction_out <= x"00000780";
when 144 => instruction_out <= x"30101831";   -- SHL R12, R12, 0x10;
when 145 => instruction_out <= x"c4100780";
when 146 => instruction_out <= x"600a0429";   -- IMAD.U16 R10, R1L, R5L, R10;
when 147 => instruction_out <= x"00028780";
when 148 => instruction_out <= x"30101a05";   -- SHL R1, R13, 0x10;
when 149 => instruction_out <= x"c4100780";
when 150 => instruction_out <= x"60060a2d";   -- IMAD.U16 R11, R2H, R3L, R11;
when 151 => instruction_out <= x"0002c780";
when 152 => instruction_out <= x"600e0c15";   -- IMAD.U16 R5, R3L, R7L, R12;
when 153 => instruction_out <= x"00030780";
when 154 => instruction_out <= x"6010181d";   -- IMAD.U16 R7, R6L, R8L, R1;
when 155 => instruction_out <= x"00004780";
when 156 => instruction_out <= x"400d1431";   -- IMUL.U16.U16 R12, R5L, R6H;
when 157 => instruction_out <= x"00000780";
when 158 => instruction_out <= x"10018005";   -- MVI R1, 0x1;
when 159 => instruction_out <= x"00000003";
when 160 => instruction_out <= x"30101621";   -- SHL R8, R11, 0x10;
when 161 => instruction_out <= x"c4100780";
when 162 => instruction_out <= x"40091c35";   -- IMUL.U16.U16 R13, R7L, R4H;
when 163 => instruction_out <= x"00000780";
when 164 => instruction_out <= x"600c162d";   -- IMAD.U16 R11, R5H, R6L, R12;
when 165 => instruction_out <= x"00030780";
when 166 => instruction_out <= x"30090205";   -- SHL R1, R1, R9;
when 167 => instruction_out <= x"c4000780";
when 168 => instruction_out <= x"6006080d";   -- IMAD.U16 R3, R2L, R3L, R8;
when 169 => instruction_out <= x"00020780";
when 170 => instruction_out <= x"60081e25";   -- IMAD.U16 R9, R7H, R4L, R13;
when 171 => instruction_out <= x"00034780";
when 172 => instruction_out <= x"30101621";   -- SHL R8, R11, 0x10;
when 173 => instruction_out <= x"c4100780";
when 174 => instruction_out <= x"301f0209";   -- SHR.S32 R2, R1, 0x1f;
when 175 => instruction_out <= x"ec100780";
when 176 => instruction_out <= x"2000140d";   -- IADD R3, R10, R3;
when 177 => instruction_out <= x"0400c780";
when 178 => instruction_out <= x"30101225";   -- SHL R9, R9, 0x10;
when 179 => instruction_out <= x"c4100780";
when 180 => instruction_out <= x"600c1415";   -- IMAD.U16 R5, R5L, R6L, R8;
when 181 => instruction_out <= x"00020780";
when 182 => instruction_out <= x"3002d7fd";   -- ISET.C1 o[0x7f], g [0xb], R2, EQ;
when 183 => instruction_out <= x"642087d8";
when 184 => instruction_out <= x"a0000001";   -- I2I.U32.U16 R0, R0L;
when 185 => instruction_out <= x"04000780";
when 186 => instruction_out <= x"60081c11";   -- IMAD.U16 R4, R7L, R4L, R9;
when 187 => instruction_out <= x"00024780";
when 188 => instruction_out <= x"20038000";   -- IADD32 R0, R0, R3;
when 189 => instruction_out <= x"20048a0c";   -- IADD32 R3, R5, R4;
when 190 => instruction_out <= x"3002d7fd";   -- ISET.C1 o[0x7f] (C1.EQ), g [0xb], R2, LT;
when 191 => instruction_out <= x"64205158";
when 192 => instruction_out <= x"2000000d";   -- IADD R3, R0, R3;
when 193 => instruction_out <= x"0400c780";
when 194 => instruction_out <= x"307ccffd";   -- ISET.S32.C0 o[0x7f], g [0x7], R124, LE;
when 195 => instruction_out <= x"6c2107c8";
when 196 => instruction_out <= x"100a2003";   -- BRA C1.NE, 0x510;
when 197 => instruction_out <= x"00001280";
when 198 => instruction_out <= x"1100ee00";   -- MOV32 R0, g [0x7];
when 199 => instruction_out <= x"10008208";   -- MOV32 R2, R1;
when 200 => instruction_out <= x"1006c003";   -- BRA C0.EQ, 0x360;
when 201 => instruction_out <= x"00000100";
when 202 => instruction_out <= x"1000f811";   -- MOV R4, R124;
when 203 => instruction_out <= x"0403c780";
when 204 => instruction_out <= x"30010001";   -- SHR.S32 R0, R0, 0x1;
when 205 => instruction_out <= x"ec100780";
when 206 => instruction_out <= x"307c01fd";   -- ISET.S32.C1 o[0x7f], R0, R124, GT;
when 207 => instruction_out <= x"6c0107d8";
when 208 => instruction_out <= x"20018811";   -- IADD32I R4, R4, 0x1;
when 209 => instruction_out <= x"00000003";
when 210 => instruction_out <= x"10067003";   -- BRA C1.NE, 0x338;
when 211 => instruction_out <= x"00001280";
when 212 => instruction_out <= x"1006d003";   -- BRA  0x368;
when 213 => instruction_out <= x"00000780";
when 214 => instruction_out <= x"1000f811";   -- MOV R4, R124;
when 215 => instruction_out <= x"0403c780";
when 216 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, LE;
when 217 => instruction_out <= x"6c00c7d8";
when 218 => instruction_out <= x"10075003";   -- BRA C1.NE, 0x3a8;
when 219 => instruction_out <= x"00001280";
when 220 => instruction_out <= x"1000f801";   -- MOV R0, R124;
when 221 => instruction_out <= x"0403c780";
when 222 => instruction_out <= x"30010409";   -- SHR.S32 R2, R2, 0x1;
when 223 => instruction_out <= x"ec100780";
when 224 => instruction_out <= x"307c05fd";   -- ISET.S32.C1 o[0x7f], R2, R124, GT;
when 225 => instruction_out <= x"6c0107d8";
when 226 => instruction_out <= x"20018001";   -- IADD32I R0, R0, 0x1;
when 227 => instruction_out <= x"00000003";
when 228 => instruction_out <= x"10070003";   -- BRA C1.NE, 0x380;
when 229 => instruction_out <= x"00001280";
when 230 => instruction_out <= x"10076003";   -- BRA  0x3b0;
when 231 => instruction_out <= x"00000780";
when 232 => instruction_out <= x"1000f801";   -- MOV R0, R124;
when 233 => instruction_out <= x"0403c780";
when 234 => instruction_out <= x"20400801";   -- IADD R0, R4, -R0;
when 235 => instruction_out <= x"04000780";
when 236 => instruction_out <= x"10018009";   -- MVI R2, 0x1;
when 237 => instruction_out <= x"00000003";
when 238 => instruction_out <= x"30000409";   -- SHL R2, R2, R0;
when 239 => instruction_out <= x"c4000780";
when 240 => instruction_out <= x"307c0401";   -- ISET.S32.C2 R0, R2, R124, GT;
when 241 => instruction_out <= x"6c0107e0";
when 242 => instruction_out <= x"a00001fd";   -- I2I.S32.S32.C1 o[0x7f], R0;
when 243 => instruction_out <= x"0c0147d8";
when 244 => instruction_out <= x"10000401";   -- MOV R0, R2;
when 245 => instruction_out <= x"0403c780";
when 246 => instruction_out <= x"10083003";   -- BRA C2.EQ, 0x418;
when 247 => instruction_out <= x"00002100";
when 248 => instruction_out <= x"1000f811";   -- MOV R4, R124;
when 249 => instruction_out <= x"0403c780";
when 250 => instruction_out <= x"30010409";   -- SHR.S32 R2, R2, 0x1;
when 251 => instruction_out <= x"ec100780";
when 252 => instruction_out <= x"307c05fd";   -- ISET.S32.C2 o[0x7f], R2, R124, GT;
when 253 => instruction_out <= x"6c0107e8";
when 254 => instruction_out <= x"20018811";   -- IADD32I R4, R4, 0x1;
when 255 => instruction_out <= x"00000003";
when 256 => instruction_out <= x"1007e003";   -- BRA C2.NE, 0x3f0;
when 257 => instruction_out <= x"00002280";
when 258 => instruction_out <= x"10084003";   -- BRA  0x420;
when 259 => instruction_out <= x"00000780";
when 260 => instruction_out <= x"1000f811";   -- MOV R4, R124;
when 261 => instruction_out <= x"0403c780";
when 262 => instruction_out <= x"203f8009";   -- IADD32I R2, R0, 0xffffffff;
when 263 => instruction_out <= x"0fffffff";
when 264 => instruction_out <= x"d0020615";   -- LOP.AND R5, R3, R2;
when 265 => instruction_out <= x"04000780";
when 266 => instruction_out <= x"400b0409";   -- IMUL.U16.U16 R2, R1L, R5H;
when 267 => instruction_out <= x"00000780";
when 268 => instruction_out <= x"600a0619";   -- IMAD.U16 R6, R1H, R5L, R2;
when 269 => instruction_out <= x"00008780";
when 270 => instruction_out <= x"203f8809";   -- IADD32I R2, R4, 0xffffffff;
when 271 => instruction_out <= x"0fffffff";
when 272 => instruction_out <= x"30100c11";   -- SHL R4, R6, 0x10;
when 273 => instruction_out <= x"c4100780";
when 274 => instruction_out <= x"30020625";   -- SHR.S32 R9, R3, R2;
when 275 => instruction_out <= x"ec000780";
when 276 => instruction_out <= x"600a0411";   -- IMAD.U16 R4, R1L, R5L, R4;
when 277 => instruction_out <= x"00010780";
when 278 => instruction_out <= x"1000ce05";   -- MOV R1, g [0x7];
when 279 => instruction_out <= x"0423c780";
when 280 => instruction_out <= x"10094003";   -- BRA C0.EQ, 0x4a0;
when 281 => instruction_out <= x"00000100";
when 282 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 283 => instruction_out <= x"0403c780";
when 284 => instruction_out <= x"30010205";   -- SHR.S32 R1, R1, 0x1;
when 285 => instruction_out <= x"ec100780";
when 286 => instruction_out <= x"307c03fd";   -- ISET.S32.C0 o[0x7f], R1, R124, GT;
when 287 => instruction_out <= x"6c0107c8";
when 288 => instruction_out <= x"20018409";   -- IADD32I R2, R2, 0x1;
when 289 => instruction_out <= x"00000003";
when 290 => instruction_out <= x"1008f003";   -- BRA C0.NE, 0x478;
when 291 => instruction_out <= x"00000280";
when 292 => instruction_out <= x"10095003";   -- BRA  0x4a8;
when 293 => instruction_out <= x"00000780";
when 294 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 295 => instruction_out <= x"0403c780";
when 296 => instruction_out <= x"1009c003";   -- BRA C1.EQ, 0x4e0;
when 297 => instruction_out <= x"00001100";
when 298 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 299 => instruction_out <= x"0403c780";
when 300 => instruction_out <= x"30010001";   -- SHR.S32 R0, R0, 0x1;
when 301 => instruction_out <= x"ec100780";
when 302 => instruction_out <= x"307c01fd";   -- ISET.S32.C0 o[0x7f], R0, R124, GT;
when 303 => instruction_out <= x"6c0107c8";
when 304 => instruction_out <= x"20018205";   -- IADD32I R1, R1, 0x1;
when 305 => instruction_out <= x"00000003";
when 306 => instruction_out <= x"10097003";   -- BRA C0.NE, 0x4b8;
when 307 => instruction_out <= x"00000280";
when 308 => instruction_out <= x"1009d003";   -- BRA  0x4e8;
when 309 => instruction_out <= x"00000780";
when 310 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 311 => instruction_out <= x"0403c780";
when 312 => instruction_out <= x"20400401";   -- IADD R0, R2, -R1;
when 313 => instruction_out <= x"04004780";
when 314 => instruction_out <= x"10018005";   -- MVI R1, 0x1;
when 315 => instruction_out <= x"00000003";
when 316 => instruction_out <= x"30000215";   -- SHL R5, R1, R0;
when 317 => instruction_out <= x"c4000780";
when 318 => instruction_out <= x"10018029";   -- MVI R10, 0x1;
when 319 => instruction_out <= x"00000003";
when 320 => instruction_out <= x"100db003";   -- BRA  0x6d8;
when 321 => instruction_out <= x"00000780";
when 322 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, LE;
when 323 => instruction_out <= x"6c00c7d8";
when 324 => instruction_out <= x"1000ce01";   -- MOV R0, g [0x7];
when 325 => instruction_out <= x"0423c780";
when 326 => instruction_out <= x"100ab003";   -- BRA C1.NE, 0x558;
when 327 => instruction_out <= x"00001280";
when 328 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 329 => instruction_out <= x"0403c780";
when 330 => instruction_out <= x"30010205";   -- SHR.S32 R1, R1, 0x1;
when 331 => instruction_out <= x"ec100780";
when 332 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, GT;
when 333 => instruction_out <= x"6c0107d8";
when 334 => instruction_out <= x"20018409";   -- IADD32I R2, R2, 0x1;
when 335 => instruction_out <= x"00000003";
when 336 => instruction_out <= x"100a6003";   -- BRA C1.NE, 0x530;
when 337 => instruction_out <= x"00001280";
when 338 => instruction_out <= x"100ac003";   -- BRA  0x560;
when 339 => instruction_out <= x"00000780";
when 340 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 341 => instruction_out <= x"0403c780";
when 342 => instruction_out <= x"100b3003";   -- BRA C0.EQ, 0x598;
when 343 => instruction_out <= x"00000100";
when 344 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 345 => instruction_out <= x"0403c780";
when 346 => instruction_out <= x"30010001";   -- SHR.S32 R0, R0, 0x1;
when 347 => instruction_out <= x"ec100780";
when 348 => instruction_out <= x"307c01fd";   -- ISET.S32.C0 o[0x7f], R0, R124, GT;
when 349 => instruction_out <= x"6c0107c8";
when 350 => instruction_out <= x"20018205";   -- IADD32I R1, R1, 0x1;
when 351 => instruction_out <= x"00000003";
when 352 => instruction_out <= x"100ae003";   -- BRA C0.NE, 0x570;
when 353 => instruction_out <= x"00000280";
when 354 => instruction_out <= x"100b4003";   -- BRA  0x5a0;
when 355 => instruction_out <= x"00000780";
when 356 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 357 => instruction_out <= x"0403c780";
when 358 => instruction_out <= x"20400401";   -- IADD R0, R2, -R1;
when 359 => instruction_out <= x"04004780";
when 360 => instruction_out <= x"10018005";   -- MVI R1, 0x1;
when 361 => instruction_out <= x"00000003";
when 362 => instruction_out <= x"30000205";   -- SHL R1, R1, R0;
when 363 => instruction_out <= x"c4000780";
when 364 => instruction_out <= x"307c0201";   -- ISET.S32.C1 R0, R1, R124, GT;
when 365 => instruction_out <= x"6c0107d0";
when 366 => instruction_out <= x"a00001fd";   -- I2I.S32.S32.C0 o[0x7f], R0;
when 367 => instruction_out <= x"0c0147c8";
when 368 => instruction_out <= x"10000201";   -- MOV R0, R1;
when 369 => instruction_out <= x"0403c780";
when 370 => instruction_out <= x"100c1003";   -- BRA C1.EQ, 0x608;
when 371 => instruction_out <= x"00001100";
when 372 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 373 => instruction_out <= x"0403c780";
when 374 => instruction_out <= x"30010205";   -- SHR.S32 R1, R1, 0x1;
when 375 => instruction_out <= x"ec100780";
when 376 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, GT;
when 377 => instruction_out <= x"6c0107d8";
when 378 => instruction_out <= x"20018409";   -- IADD32I R2, R2, 0x1;
when 379 => instruction_out <= x"00000003";
when 380 => instruction_out <= x"100bc003";   -- BRA C1.NE, 0x5e0;
when 381 => instruction_out <= x"00001280";
when 382 => instruction_out <= x"100c2003";   -- BRA  0x610;
when 383 => instruction_out <= x"00000780";
when 384 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 385 => instruction_out <= x"0403c780";
when 386 => instruction_out <= x"203f8405";   -- IADD32I R1, R2, 0xffffffff;
when 387 => instruction_out <= x"0fffffff";
when 388 => instruction_out <= x"307ccdfd";   -- ISET.S32.C0 o[0x7f], g [0x6], R124, LE;
when 389 => instruction_out <= x"6c20c7d8";
when 390 => instruction_out <= x"30010625";   -- SHL R9, R3, R1;
when 391 => instruction_out <= x"c4000780";
when 392 => instruction_out <= x"1000cc05";   -- MOV R1, g [0x6];
when 393 => instruction_out <= x"0423c780";
when 394 => instruction_out <= x"100cd003";   -- BRA C1.NE, 0x668;
when 395 => instruction_out <= x"00001280";
when 396 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 397 => instruction_out <= x"0403c780";
when 398 => instruction_out <= x"30010205";   -- SHR.S32 R1, R1, 0x1;
when 399 => instruction_out <= x"ec100780";
when 400 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, GT;
when 401 => instruction_out <= x"6c0107d8";
when 402 => instruction_out <= x"20018409";   -- IADD32I R2, R2, 0x1;
when 403 => instruction_out <= x"00000003";
when 404 => instruction_out <= x"100c8003";   -- BRA C1.NE, 0x640;
when 405 => instruction_out <= x"00001280";
when 406 => instruction_out <= x"100ce003";   -- BRA  0x670;
when 407 => instruction_out <= x"00000780";
when 408 => instruction_out <= x"1000f809";   -- MOV R2, R124;
when 409 => instruction_out <= x"0403c780";
when 410 => instruction_out <= x"100d5003";   -- BRA C0.EQ, 0x6a8;
when 411 => instruction_out <= x"00000100";
when 412 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 413 => instruction_out <= x"0403c780";
when 414 => instruction_out <= x"30010001";   -- SHR.S32 R0, R0, 0x1;
when 415 => instruction_out <= x"ec100780";
when 416 => instruction_out <= x"307c01fd";   -- ISET.S32.C0 o[0x7f], R0, R124, GT;
when 417 => instruction_out <= x"6c0107c8";
when 418 => instruction_out <= x"20018205";   -- IADD32I R1, R1, 0x1;
when 419 => instruction_out <= x"00000003";
when 420 => instruction_out <= x"100d0003";   -- BRA C0.NE, 0x680;
when 421 => instruction_out <= x"00000280";
when 422 => instruction_out <= x"100d6003";   -- BRA  0x6b0;
when 423 => instruction_out <= x"00000780";
when 424 => instruction_out <= x"1000f805";   -- MOV R1, R124;
when 425 => instruction_out <= x"0403c780";
when 426 => instruction_out <= x"20400401";   -- IADD R0, R2, -R1;
when 427 => instruction_out <= x"04004780";
when 428 => instruction_out <= x"10018005";   -- MVI R1, 0x1;
when 429 => instruction_out <= x"00000003";
when 430 => instruction_out <= x"30000229";   -- SHL R10, R1, R0;
when 431 => instruction_out <= x"c4000780";
when 432 => instruction_out <= x"1000ce15";   -- MOV R5, g [0x7];
when 433 => instruction_out <= x"0423c780";
when 434 => instruction_out <= x"1000f811";   -- MOV R4, R124;
when 435 => instruction_out <= x"0403c780";
when 436 => instruction_out <= x"307c1401";   -- ISET.S32.C1 R0, R10, R124, GT;
when 437 => instruction_out <= x"6c0107d0";
when 438 => instruction_out <= x"a00001fd";   -- I2I.S32.S32.C0 o[0x7f], R0;
when 439 => instruction_out <= x"0c0147c8";
when 440 => instruction_out <= x"10109003";   -- BRA C1.EQ, 0x848;
when 441 => instruction_out <= x"00001100";
when 442 => instruction_out <= x"307c0bfd";   -- ISET.S32.C1 o[0x7f], R5, R124, GT;
when 443 => instruction_out <= x"6c0107d8";
when 444 => instruction_out <= x"1000f821";   -- MOV R8, R124;
when 445 => instruction_out <= x"0403c780";
when 446 => instruction_out <= x"10106003";   -- BRA C1.EQ, 0x830;
when 447 => instruction_out <= x"00001100";
when 448 => instruction_out <= x"20001201";   -- IADD R0, R9, R8;
when 449 => instruction_out <= x"04020780";
when 450 => instruction_out <= x"3004002d";   -- SHL R11, R0, 0x4;
when 451 => instruction_out <= x"c4100780";
when 452 => instruction_out <= x"30050001";   -- SHL R0, R0, 0x5;
when 453 => instruction_out <= x"c4100780";
when 454 => instruction_out <= x"30010805";   -- SHL R1, R4, 0x1;
when 455 => instruction_out <= x"c4100780";
when 456 => instruction_out <= x"200b8000";   -- IADD32 R0, R0, R11;
when 457 => instruction_out <= x"20048204";   -- IADD32 R1, R1, R4;
when 458 => instruction_out <= x"2100e800";   -- IADD32 R0, g [0x4], R0;
when 459 => instruction_out <= x"20018030";   -- IADD32 R12, R0, R1;
when 460 => instruction_out <= x"a0105003";   -- SSY 0x828;
when 461 => instruction_out <= x"00000000";
when 462 => instruction_out <= x"10008804";   -- MOV32 R1, R4;
when 463 => instruction_out <= x"20058834";   -- IADD32 R13, R4, R5;
when 464 => instruction_out <= x"10000809";   -- MOV R2, R4;
when 465 => instruction_out <= x"0403c780";
when 466 => instruction_out <= x"d00e1801";   -- GLD.U8 R0, global14[R12];
when 467 => instruction_out <= x"80000780";
when 468 => instruction_out <= x"2001980d";   -- IADD32I R3, R12, 0x1;
when 469 => instruction_out <= x"00000003";
when 470 => instruction_out <= x"d00e060d";   -- GLD.U8 R3, global14[R3];
when 471 => instruction_out <= x"80000780";
when 472 => instruction_out <= x"20029819";   -- IADD32I R6, R12, 0x2;
when 473 => instruction_out <= x"00000003";
when 474 => instruction_out <= x"d00e0c1d";   -- GLD.U8 R7, global14[R6];
when 475 => instruction_out <= x"80000780";
when 476 => instruction_out <= x"10058019";   -- MVI R6, 0x9645;
when 477 => instruction_out <= x"00000967";
when 478 => instruction_out <= x"40061a39";   -- IMUL.U16.U16 R14, R6H, R3L;
when 479 => instruction_out <= x"00000780";
when 480 => instruction_out <= x"30101c39";   -- SHL R14, R14, 0x10;
when 481 => instruction_out <= x"c4100780";
when 482 => instruction_out <= x"40048101";   -- IMUL32I.S16.S16 R0, R0L, 0x4c84;
when 483 => instruction_out <= x"000004cb";
when 484 => instruction_out <= x"6006180d";   -- IMAD.U16 R3, R6L, R3L, R14;
when 485 => instruction_out <= x"00038780";
when 486 => instruction_out <= x"30100001";   -- SHR.S32 R0, R0, 0x10;
when 487 => instruction_out <= x"ec100780";
when 488 => instruction_out <= x"3010060d";   -- SHR.S32 R3, R3, 0x10;
when 489 => instruction_out <= x"ec100780";
when 490 => instruction_out <= x"401f9d19";   -- IMUL32I.S16.S16 R6, R7L, 0x12df;
when 491 => instruction_out <= x"0000012f";
when 492 => instruction_out <= x"20000001";   -- IADD R0, R0, R3;
when 493 => instruction_out <= x"0400c780";
when 494 => instruction_out <= x"30100c0d";   -- SHR.S32 R3, R6, 0x10;
when 495 => instruction_out <= x"ec100780";
when 496 => instruction_out <= x"20000001";   -- IADD R0, R0, R3;
when 497 => instruction_out <= x"0400c780";
when 498 => instruction_out <= x"a0000001";   -- I2I.S32.S16 R0, R0L;
when 499 => instruction_out <= x"0c010780";
when 500 => instruction_out <= x"20018205";   -- IADD32I R1, R1, 0x1;
when 501 => instruction_out <= x"00000003";
when 502 => instruction_out <= x"2000040d";   -- IADD R3, R2, R11;
when 503 => instruction_out <= x"0402c780";
when 504 => instruction_out <= x"308101fd";   -- ISET.S32.C2 o[0x7f], R0, c[0x1][0x1], GT;
when 505 => instruction_out <= x"6c4107e8";
when 506 => instruction_out <= x"10000201";   -- MVC R0 (C2.NE), c[0x1] [0x1];
when 507 => instruction_out <= x"2440e280";
when 508 => instruction_out <= x"300d03fd";   -- ISET.S32.C2 o[0x7f], R1, R13, NE;
when 509 => instruction_out <= x"6c0147e8";
when 510 => instruction_out <= x"2100060d";   -- IADD R3, R3, c[0xe][0x0];
when 511 => instruction_out <= x"07800780";
when 512 => instruction_out <= x"d00e0601";   -- GST.U8 global14[R3], R0;
when 513 => instruction_out <= x"a0000780";
when 514 => instruction_out <= x"20018409";   -- IADD32I R2, R2, 0x1;
when 515 => instruction_out <= x"00000003";
when 516 => instruction_out <= x"20039831";   -- IADD32I R12, R12, 0x3;
when 517 => instruction_out <= x"00000003";
when 518 => instruction_out <= x"100ea003";   -- BRA C2.NE, 0x750;
when 519 => instruction_out <= x"00002280";
when 520 => instruction_out <= x"f0000001";   -- NOP.S;
when 521 => instruction_out <= x"e0000002";
when 522 => instruction_out <= x"20019021";   -- IADD32I R8, R8, 0x1;
when 523 => instruction_out <= x"00000003";
when 524 => instruction_out <= x"300a11fd";   -- ISET.S32.C2 o[0x7f], R8, R10, NE;
when 525 => instruction_out <= x"6c0147e8";
when 526 => instruction_out <= x"100e0003";   -- BRA C2.NE, 0x700;
when 527 => instruction_out <= x"00002280";
when 528 => instruction_out <= x"30000003";   -- RET C0.EQ;
when 529 => instruction_out <= x"00000100";
when 530 => instruction_out <= x"307c0bfd";   -- ISET.S32.C0 o[0x7f], R5, R124, GT;
when 531 => instruction_out <= x"6c0107c8";
when 532 => instruction_out <= x"1000f82d";   -- MOV R11, R124;
when 533 => instruction_out <= x"0403c780";
when 534 => instruction_out <= x"10169003";   -- BRA C0.EQ, 0xb48;
when 535 => instruction_out <= x"00000100";
when 536 => instruction_out <= x"20001201";   -- IADD R0, R9, R11;
when 537 => instruction_out <= x"0402c780";
when 538 => instruction_out <= x"21000009";   -- IADD.C1 R2, R0, c[0x1][0x2];
when 539 => instruction_out <= x"044087d0";
when 540 => instruction_out <= x"301f0005";   -- SHR.S32 R1, R0, 0x1f;
when 541 => instruction_out <= x"ec100780";
when 542 => instruction_out <= x"3140d21d";   -- IADD.CARRY2 R7, g [0x9], c[0x1][0x3];
when 543 => instruction_out <= x"0460e780";
when 544 => instruction_out <= x"3040020d";   -- IADD.CARRY1 R3, R1, R124;
when 545 => instruction_out <= x"041f1780";
when 546 => instruction_out <= x"30060431";   -- ISET R12, R2, R6, LE;
when 547 => instruction_out <= x"6400c780";
when 548 => instruction_out <= x"203f9205";   -- IADD32I R1, R9, 0xffffffff;
when 549 => instruction_out <= x"0fffffff";
when 550 => instruction_out <= x"30070621";   -- ISET R8, R3, R7, EQ;
when 551 => instruction_out <= x"64008780";
when 552 => instruction_out <= x"30070609";   -- ISET R2, R3, R7, LT;
when 553 => instruction_out <= x"64004780";
when 554 => instruction_out <= x"20001605";   -- IADD R1, R11, R1;
when 555 => instruction_out <= x"04004780";
when 556 => instruction_out <= x"d00c100d";   -- LOP.AND R3, R8, R12;
when 557 => instruction_out <= x"04000780";
when 558 => instruction_out <= x"3140d61d";   -- IADD.CARRY1 R7, g [0xb], c[0x1][0x3];
when 559 => instruction_out <= x"0460d780";
when 560 => instruction_out <= x"307c03fd";   -- ISET.S32.C1 o[0x7f], R1, R124, GE;
when 561 => instruction_out <= x"6c0187d8";
when 562 => instruction_out <= x"d00305fd";   -- LOP.OR.C2 o[0x7f], R2, R3;
when 563 => instruction_out <= x"040047e8";
when 564 => instruction_out <= x"a0168003";   -- SSY 0xb40;
when 565 => instruction_out <= x"00000000";
when 566 => instruction_out <= x"30040039";   -- SHL R14, R0, 0x4;
when 567 => instruction_out <= x"c4100780";
when 568 => instruction_out <= x"1000883c";   -- MOV32 R15, R4;
when 569 => instruction_out <= x"20058840";   -- IADD32 R16, R4, R5;
when 570 => instruction_out <= x"203f8845";   -- IADD32I R17, R4, 0xffffffff;
when 571 => instruction_out <= x"0fffffff";
when 572 => instruction_out <= x"210eea00";   -- IADD32 R0, g [0x5], R14;
when 573 => instruction_out <= x"10008808";   -- MOV32 R2, R4;
when 574 => instruction_out <= x"301f080d";   -- SHR.S32 R3, R4, 0x1f;
when 575 => instruction_out <= x"ec100780";
when 576 => instruction_out <= x"21001c35";   -- IADD R13, R14, c[0xe][0x0];
when 577 => instruction_out <= x"07800780";
when 578 => instruction_out <= x"20000831";   -- IADD R12, R4, R0;
when 579 => instruction_out <= x"04000780";
when 580 => instruction_out <= x"20000401";   -- IADD R0, R2, R13;
when 581 => instruction_out <= x"04034780";
when 582 => instruction_out <= x"d00e0001";   -- GLD.U8 R0, global14[R0];
when 583 => instruction_out <= x"80000780";
when 584 => instruction_out <= x"403c8105";   -- IMUL32I.S16.S16 R1, R0L, 0xfffffffc;
when 585 => instruction_out <= x"0fffffff";
when 586 => instruction_out <= x"21000401";   -- IADD.C3 R0, R2, c[0x1][0x2];
when 587 => instruction_out <= x"044087f0";
when 588 => instruction_out <= x"30400621";   -- IADD.CARRY3 R8, R3, R124;
when 589 => instruction_out <= x"041f3780";
when 590 => instruction_out <= x"300711fd";   -- ISET.C3 o[0x7f], R8, R7, EQ;
when 591 => instruction_out <= x"640087f8";
when 592 => instruction_out <= x"300601fd";   -- ISET.C3 o[0x7f] (C3.NE), R0, R6, GT;
when 593 => instruction_out <= x"640132f8";
when 594 => instruction_out <= x"300711fd";   -- ISET.C3 o[0x7f] (C3.EQ), R8, R7, GT;
when 595 => instruction_out <= x"64013178";
when 596 => instruction_out <= x"a000040d";   -- I2I.S32.S16 R3, R1L;
when 597 => instruction_out <= x"0c010780";
when 598 => instruction_out <= x"a0138003";   -- SSY 0x9c0;
when 599 => instruction_out <= x"00000000";
when 600 => instruction_out <= x"10001005";   -- MOV R1, R8;
when 601 => instruction_out <= x"0403c780";
when 602 => instruction_out <= x"10138003";   -- BRA C3.NE, 0x9c0;
when 603 => instruction_out <= x"00003280";
when 604 => instruction_out <= x"20000421";   -- IADD R8, R2, R14;
when 605 => instruction_out <= x"04038780";
when 606 => instruction_out <= x"21001021";   -- IADD R8, R8, c[0xe][0x0];
when 607 => instruction_out <= x"07800780";
when 608 => instruction_out <= x"20019021";   -- IADD32I R8, R8, 0x1;
when 609 => instruction_out <= x"00000003";
when 610 => instruction_out <= x"d00e1021";   -- GLD.U8 R8, global14[R8];
when 611 => instruction_out <= x"80000780";
when 612 => instruction_out <= x"a0002021";   -- I2I.U32.U16.BEXT R8, R8L;
when 613 => instruction_out <= x"04008780";
when 614 => instruction_out <= x"2000060d";   -- IADD R3, R3, R8;
when 615 => instruction_out <= x"04020780";
when 616 => instruction_out <= x"a0000c0d";   -- I2I.S32.S16 R3, R3L;
when 617 => instruction_out <= x"0c010780";
when 618 => instruction_out <= x"f0000001";   -- NOP.S;
when 619 => instruction_out <= x"e0000002";
when 620 => instruction_out <= x"a0142003";   -- SSY 0xa10;
when 621 => instruction_out <= x"00000000";
when 622 => instruction_out <= x"10142003";   -- BRA C2.EQ, 0xa10;
when 623 => instruction_out <= x"00002100";
when 624 => instruction_out <= x"20000421";   -- IADD R8, R2, R14;
when 625 => instruction_out <= x"04038780";
when 626 => instruction_out <= x"21001021";   -- IADD R8, R8, c[0xe][0x0];
when 627 => instruction_out <= x"07800780";
when 628 => instruction_out <= x"20109021";   -- IADD32I R8, R8, 0x10;
when 629 => instruction_out <= x"00000003";
when 630 => instruction_out <= x"d00e1021";   -- GLD.U8 R8, global14[R8];
when 631 => instruction_out <= x"80000780";
when 632 => instruction_out <= x"a0002021";   -- I2I.U32.U16.BEXT R8, R8L;
when 633 => instruction_out <= x"04008780";
when 634 => instruction_out <= x"2000060d";   -- IADD R3, R3, R8;
when 635 => instruction_out <= x"04020780";
when 636 => instruction_out <= x"a0000c0d";   -- I2I.S32.S16 R3, R3L;
when 637 => instruction_out <= x"0c010780";
when 638 => instruction_out <= x"f0000001";   -- NOP.S;
when 639 => instruction_out <= x"e0000002";
when 640 => instruction_out <= x"a014d003";   -- SSY 0xa68;
when 641 => instruction_out <= x"00000000";
when 642 => instruction_out <= x"307c23fd";   -- ISET.S32.C3 o[0x7f], R17, R124, LT;
when 643 => instruction_out <= x"6c0047f8";
when 644 => instruction_out <= x"1014d003";   -- BRA C3.NE, 0xa68;
when 645 => instruction_out <= x"00003280";
when 646 => instruction_out <= x"20000421";   -- IADD R8, R2, R14;
when 647 => instruction_out <= x"04038780";
when 648 => instruction_out <= x"21001021";   -- IADD R8, R8, c[0xe][0x0];
when 649 => instruction_out <= x"07800780";
when 650 => instruction_out <= x"203f9021";   -- IADD32I R8, R8, 0xffffffff;
when 651 => instruction_out <= x"0fffffff";
when 652 => instruction_out <= x"d00e1021";   -- GLD.U8 R8, global14[R8];
when 653 => instruction_out <= x"80000780";
when 654 => instruction_out <= x"a0002021";   -- I2I.U32.U16.BEXT R8, R8L;
when 655 => instruction_out <= x"04008780";
when 656 => instruction_out <= x"2000060d";   -- IADD R3, R3, R8;
when 657 => instruction_out <= x"04020780";
when 658 => instruction_out <= x"a0000c0d";   -- I2I.S32.S16 R3, R3L;
when 659 => instruction_out <= x"0c010780";
when 660 => instruction_out <= x"f0000001";   -- NOP.S;
when 661 => instruction_out <= x"e0000002";
when 662 => instruction_out <= x"a0157003";   -- SSY 0xab8;
when 663 => instruction_out <= x"00000000";
when 664 => instruction_out <= x"10157003";   -- BRA C1.EQ, 0xab8;
when 665 => instruction_out <= x"00001100";
when 666 => instruction_out <= x"20000409";   -- IADD R2, R2, R14;
when 667 => instruction_out <= x"04038780";
when 668 => instruction_out <= x"21000409";   -- IADD R2, R2, c[0xe][0x0];
when 669 => instruction_out <= x"07800780";
when 670 => instruction_out <= x"20308409";   -- IADD32I R2, R2, 0xfffffff0;
when 671 => instruction_out <= x"0fffffff";
when 672 => instruction_out <= x"d00e0409";   -- GLD.U8 R2, global14[R2];
when 673 => instruction_out <= x"80000780";
when 674 => instruction_out <= x"a0000809";   -- I2I.U32.U16.BEXT R2, R2L;
when 675 => instruction_out <= x"04008780";
when 676 => instruction_out <= x"20000609";   -- IADD R2, R3, R2;
when 677 => instruction_out <= x"04008780";
when 678 => instruction_out <= x"a000080d";   -- I2I.S32.S16 R3, R2L;
when 679 => instruction_out <= x"0c010780";
when 680 => instruction_out <= x"f0000001";   -- NOP.S;
when 681 => instruction_out <= x"e0000002";
when 682 => instruction_out <= x"a015f003";   -- SSY 0xaf8;
when 683 => instruction_out <= x"00000000";
when 684 => instruction_out <= x"307c07fd";   -- ISET.S32.C3 o[0x7f], R3, R124, GE;
when 685 => instruction_out <= x"6c0187f8";
when 686 => instruction_out <= x"1015d003";   -- BRA C3.NE, 0xae8;
when 687 => instruction_out <= x"00003280";
when 688 => instruction_out <= x"1000f80d";   -- MOV R3, R124;
when 689 => instruction_out <= x"0403c780";
when 690 => instruction_out <= x"1015f003";   -- BRA  0xaf8;
when 691 => instruction_out <= x"00000780";
when 692 => instruction_out <= x"308107fd";   -- ISET.S32.C3 o[0x7f], R3, c[0x1][0x1], LE;
when 693 => instruction_out <= x"6c40c7f8";
when 694 => instruction_out <= x"1000020d";   -- MVC R3 (C3.EQU), c[0x1] [0x1];
when 695 => instruction_out <= x"2440f500";
when 696 => instruction_out <= x"f0000001";   -- NOP.S;
when 697 => instruction_out <= x"e0000002";
when 698 => instruction_out <= x"10000c11";   -- MOV.U16 R2L, R3L;
when 699 => instruction_out <= x"0003c780";
when 700 => instruction_out <= x"d00e1809";   -- GST.U8 global14[R12], R2;
when 701 => instruction_out <= x"a0000780";
when 702 => instruction_out <= x"2001a245";   -- IADD32I R17, R17, 0x1;
when 703 => instruction_out <= x"00000003";
when 704 => instruction_out <= x"20019e3d";   -- IADD32I R15, R15, 0x1;
when 705 => instruction_out <= x"00000003";
when 706 => instruction_out <= x"20019831";   -- IADD32I R12, R12, 0x1;
when 707 => instruction_out <= x"00000003";
when 708 => instruction_out <= x"1000820c";   -- MOV32 R3, R1;
when 709 => instruction_out <= x"10008008";   -- MOV32 R2, R0;
when 710 => instruction_out <= x"30101ffd";   -- ISET.S32.C3 o[0x7f], R15, R16, NE;
when 711 => instruction_out <= x"6c0147f8";
when 712 => instruction_out <= x"10125003";   -- BRA C3.NE, 0x928;
when 713 => instruction_out <= x"00003280";
when 714 => instruction_out <= x"f0000001";   -- NOP.S;
when 715 => instruction_out <= x"e0000002";
when 716 => instruction_out <= x"2001962d";   -- IADD32I R11, R11, 0x1;
when 717 => instruction_out <= x"00000003";
when 718 => instruction_out <= x"300a17fd";   -- ISET.S32.C1 o[0x7f], R11, R10, NE;
when 719 => instruction_out <= x"6c0147d8";
when 720 => instruction_out <= x"1010c003";   -- BRA C1.NE, 0x860;
when 721 => instruction_out <= x"00001280";
when 722 => instruction_out <= x"f0000001";   -- NOP;
when 723 => instruction_out <= x"e0000001";
when 724 => instruction_out <= x"30000003";   -- RET
when 725 => instruction_out <= x"00000780";

			when others => null;
		end case;
	end process;

end arch;
