library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_cos is
	generic(
		word_bits	:natural:=18;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_cos is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"000000000000000000",
		"000000111111111111",
		"000001111111111110",
		"000010111111111011",
		"000011111111110101",
		"000100111111101011",
		"000101111111011100",
		"000110111111000111",
		"000111111110101011",
		"001000111110000111",
		"001001111101011010",
		"001010111100100011",
		"001011111011100001",
		"001100111010010011",
		"001101111000111001",
		"001110110111010000",
		"001111110101011000",
		"010000110011010001",
		"010001110000111001",
		"010010101110001111",
		"010011101011010011",
		"010100101000000010",
		"010101100100011101",
		"010110100000100011",
		"010111011100010010",
		"011000010111101001",
		"011001010010101001",
		"011010001101001111",
		"011011000111011010",
		"011100000001001011",
		"011100111010011111",
		"011101110011010111",
		"011110101011110001",
		"011111100011101100",
		"100000011011001000",
		"100001010010000011",
		"100010001000011101",
		"100010111110010101",
		"100011110011101001",
		"100100101000011010",
		"100101011100100111",
		"100110010000001110",
		"100111000011001110",
		"100111110101101000",
		"101000100111011010",
		"101001011000100011",
		"101010001001000011",
		"101010111000111000",
		"101011101000000011",
		"101100010110100010",
		"101101000100010101",
		"101101110001011011",
		"101110011101110011",
		"101111001001011100",
		"101111110100010111",
		"110000011110100001",
		"110001000111111011",
		"110001110000100100",
		"110010011000011011",
		"110010111111100000",
		"110011100101110010",
		"110100001011010000",
		"110100101111111010",
		"110101010011101111"
	);
begin
	data <= "10"&rom(to_integer(unsigned(addr)));
end architecture;