library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_ln2 is
	generic(
		word_bits	:natural:=27;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_ln2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"000000000000000000000000000",
		"000000101101111111001010000",
		"000001011011100111100101100",
		"000010001000111001101001000",
		"000010110101110101101001110",
		"000011100010011011111101010",
		"000100001110101100111000100",
		"000100111010101000101111110",
		"000101100110001111110111000",
		"000110010001100010100001100",
		"000110111100100001000010010",
		"000111100111001011101100000",
		"001000010001100010110001000",
		"001000111011100110100011010",
		"001001100101010111010011110",
		"001010001110110101010100000",
		"001010111000000000110100100",
		"001011100000111010000101100",
		"001100001001100001010111100",
		"001100110001110110111010000",
		"001101011001111010111100010",
		"001110000001101101101101100",
		"001110101001001111011100100",
		"001111010000100000010111110",
		"001111110111100000101101100",
		"010000011110010000101011100",
		"010001000100110000011111010",
		"010001101011000000010110110",
		"010010010001000000011110100",
		"010010110110110001000100000",
		"010011011100010010010011010",
		"010100000001100100011000110",
		"010100100110100111100001000",
		"010101001011011011111000000",
		"010101110000000001101000110",
		"010110010100011000111111100",
		"010110111000100010000111010",
		"010111011100011101001010110",
		"011000000000001010010101100",
		"011000100011101001110001110",
		"011001000110111011101010000",
		"011001101010000000001000110",
		"011010001100110111011000000",
		"011010101111100001100001110",
		"011011010001111110101111110",
		"011011110100001111001011100",
		"011100010110010010111110110",
		"011100111000001010010010010",
		"011101011001110101001111100",
		"011101111011010011111111010",
		"011110011100100110101010100",
		"011110111101101101011001110",
		"011111011110101000010101100",
		"011111111111010111100110010",
		"100000011111111011010100010",
		"100001000000010011100111100",
		"100001100000100000101000000",
		"100010000000100010011101100",
		"100010100000011001001111110",
		"100011000000000101000110100",
		"100011011111100110001000110",
		"100011111110111100011110100",
		"100100011110001000001110100",
		"100100111101001001100000000",
		"100101011100000000011010010",
		"100101111010101101000011100",
		"100110011001001111100011010",
		"100110110111100111111111110",
		"100111010101110110011111110",
		"100111110011111011001001110",
		"101000010001110110000011110",
		"101000101111100111010100110",
		"101001001101001111000010010",
		"101001101010101101010010110",
		"101010001000000010001100010",
		"101010100101001101110100010",
		"101011000010010000010001000",
		"101011011111001001101000010",
		"101011111011111001111111100",
		"101100011000100001011100100",
		"101100110101000000000100010",
		"101101010001010101111100110",
		"101101101101100011001011010",
		"101110001001100111110100110",
		"101110100101100011111110100",
		"101111000001010111101110000",
		"101111011101000011000111110",
		"101111111000100110010001000",
		"110000010100000001001110100",
		"110000101111010100000101100",
		"110001001010011110111010010",
		"110001100101100001110001110",
		"110010000000011100110000100",
		"110010011011001111111011010",
		"110010110101111011010110100",
		"110011010000011111000110100",
		"110011101010111011001111110",
		"110100000101001111110110110",
		"110100011111011100111111100",
		"110100111001100010101110100",
		"110101010011100001000111100",
		"110101101101011000001111000",
		"110110000111001000001001000",
		"110110100000110000111001100",
		"110110111010010010100100100",
		"110111010011101101001101100",
		"110111101101000000111000110",
		"111000000110001101101010000",
		"111000011111010011100101000",
		"111000111000010010101101010",
		"111001010001001011000110110",
		"111001101001111100110101000",
		"111010000010100111111011010",
		"111010011011001100011101100",
		"111010110011101010011111000",
		"111011001100000010000011000",
		"111011100100010011001101010",
		"111011111100011110000001000",
		"111100010100100010100001010",
		"111100101100100000110001110",
		"111101000100011000110101100",
		"111101011100001010101111110",
		"111101110011110110100011100",
		"111110001011011100010100000",
		"111110100010111100000100010",
		"111110111010010101110111100",
		"111111010001101001110000100",
		"111111101000110111110010010"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)));
end architecture;