library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C2_reci_sqrt_2_4 is
	generic(
		word_bits	:natural:=12;
		bus_bits	:natural:=14;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C2_reci_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"100001100000",
		"100000111000",
		"100000010000",
		"011111101000",
		"011111001000",
		"011110100000",
		"011101111000",
		"011101011000",
		"011100111000",
		"011100011000",
		"011011110000",
		"011011010000",
		"011010111000",
		"011010011000",
		"011001111000",
		"011001100000",
		"011001000000",
		"011000101000",
		"011000001000",
		"010111110000",
		"010111011000",
		"010111000000",
		"010110101000",
		"010110010000",
		"010101111000",
		"010101100000",
		"010101001000",
		"010100110000",
		"010100100000",
		"010100001000",
		"010011111000",
		"010011100000",
		"010011010000",
		"010010111000",
		"010010101000",
		"010010011000",
		"010010001000",
		"010001110000",
		"010001100000",
		"010001010000",
		"010001000000",
		"010000110000",
		"010000100000",
		"010000010000",
		"010000000000",
		"001111110000",
		"001111101000",
		"001111011000",
		"001111001000",
		"001110111000",
		"001110110000",
		"001110100000",
		"001110010000",
		"001110001000",
		"001101111000",
		"001101110000",
		"001101100000",
		"001101011000",
		"001101001000",
		"001101000000",
		"001100111000",
		"001100101000",
		"001100100000",
		"001100011000",
		"001100001000",
		"001100000000",
		"001011111000",
		"001011110000",
		"001011100000",
		"001011011000",
		"001011010000",
		"001011001000",
		"001011000000",
		"001010111000",
		"001010110000",
		"001010101000",
		"001010100000",
		"001010011000",
		"001010010000",
		"001010001000",
		"001010000000",
		"001001111000",
		"001001110000",
		"001001101000",
		"001001100000",
		"001001011000",
		"001001010000",
		"001001001000",
		"001001000000",
		"001001000000",
		"001000111000",
		"001000110000",
		"001000101000",
		"001000100000",
		"001000100000",
		"001000011000",
		"001000010000",
		"001000001000",
		"001000001000",
		"001000000000",
		"000111111000",
		"000111111000",
		"000111110000",
		"000111101000",
		"000111101000",
		"000111100000",
		"000111011000",
		"000111011000",
		"000111010000",
		"000111001000",
		"000111001000",
		"000111000000",
		"000111000000",
		"000110111000",
		"000110110000",
		"000110110000",
		"000110101000",
		"000110101000",
		"000110100000",
		"000110100000",
		"000110011000",
		"000110011000",
		"000110010000",
		"000110010000",
		"000110001000",
		"000110001000",
		"000110000000",
		"000110000000"
	);
begin
	data <= "00"&rom(to_integer(unsigned(addr)));
end architecture;