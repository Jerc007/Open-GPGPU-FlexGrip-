library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_reci_sqrt_1_2 is
	generic(
		word_bits	:natural:=17;
		bus_bits	:natural:=20;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_reci_sqrt_1_2 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"11111111111111100",
		"11111101000001100",
		"11111010000111000",
		"11110111010000000",
		"11110100011100100",
		"11110001101100100",
		"11101110111111100",
		"11101100010110000",
		"11101001101111100",
		"11100111001100000",
		"11100100101011100",
		"11100010001101100",
		"11011111110011000",
		"11011101011010100",
		"11011011000101100",
		"11011000110010100",
		"11010110100010000",
		"11010100010100100",
		"11010010001001000",
		"11010000000000000",
		"11001101111001100",
		"11001011110101000",
		"11001001110010100",
		"11000111110010100",
		"11000101110100100",
		"11000011111000100",
		"11000001111111000",
		"11000000000111000",
		"10111110010001000",
		"10111100011100100",
		"10111010101010100",
		"10111000111010000",
		"10110111001011000",
		"10110101011110000",
		"10110011110010100",
		"10110010001001000",
		"10110000100001000",
		"10101110111010000",
		"10101101010101000",
		"10101011110001100",
		"10101010001111100",
		"10101000101111000",
		"10100111010000000",
		"10100101110010000",
		"10100100010110000",
		"10100010111011000",
		"10100001100001000",
		"10100000001000100",
		"10011110110001100",
		"10011101011011100",
		"10011100000110100",
		"10011010110011000",
		"10011001100000100",
		"10011000001111000",
		"10010110111111000",
		"10010101110000000",
		"10010100100010000",
		"10010011010101000",
		"10010010001001000",
		"10010000111110000",
		"10001111110100000",
		"10001110101011000",
		"10001101100011000",
		"10001100011100000",
		"10001011010110000",
		"10001010010001000",
		"10001001001100100",
		"10001000001001000",
		"10000111000110100",
		"10000110000100100",
		"10000101000011100",
		"10000100000011100",
		"10000011000100100",
		"10000010000110000",
		"10000001001000000",
		"10000000001011000",
		"01111111001111000",
		"01111110010011100",
		"01111101011000100",
		"01111100011110100",
		"01111011100101000",
		"01111010101100100",
		"01111001110100100",
		"01111000111101000",
		"01111000000110000",
		"01110111010000000",
		"01110110011010100",
		"01110101100110000",
		"01110100110001100",
		"01110011111110000",
		"01110011001011000",
		"01110010011000100",
		"01110001100111000",
		"01110000110101100",
		"01110000000101000",
		"01101111010100100",
		"01101110100101000",
		"01101101110110000",
		"01101101000111000",
		"01101100011001000",
		"01101011101011100",
		"01101010111110100",
		"01101010010010000",
		"01101001100101100",
		"01101000111010000",
		"01101000001111000",
		"01100111100100000",
		"01100110111010000",
		"01100110010000000",
		"01100101100110100",
		"01100100111101100",
		"01100100010101000",
		"01100011101101000",
		"01100011000101100",
		"01100010011110000",
		"01100001110111100",
		"01100001010001000",
		"01100000101011000",
		"01100000000101000",
		"01011111100000000",
		"01011110111011000",
		"01011110010110100",
		"01011101110010000",
		"01011101001110100",
		"01011100101011000",
		"01011100000111100",
		"01011011100101000",
		"01011011000010100"
	);
begin
	data <= "100"&rom(to_integer(unsigned(addr)));
end architecture;