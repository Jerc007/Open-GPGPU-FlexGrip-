
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TP_instructions is
	port(
		instruction_pointer_in : in  integer;
		num_instructions_out   : out integer;
		instruction_out        : out std_logic_vector(31 downto 0)
	);
end TP_instructions;

architecture arch of TP_instructions is
	constant TP_INSTRUCTIONS : integer := 714;

begin
	num_instructions_out <= TP_INSTRUCTIONS;

	process(instruction_pointer_in)
	begin
		case instruction_pointer_in is
			when 0 => instruction_out <= x"a000440d";
when 1 => instruction_out <= x"04200780";
when 2 => instruction_out <= x"a0004219";
when 3 => instruction_out <= x"04200780";
when 4 => instruction_out <= x"400d0c05";
when 5 => instruction_out <= x"00000780";
when 6 => instruction_out <= x"600c0e05";
when 7 => instruction_out <= x"00004780";
when 8 => instruction_out <= x"30100205";
when 9 => instruction_out <= x"c4100780";
when 10 => instruction_out <= x"a0004615";
when 11 => instruction_out <= x"04200780";
when 12 => instruction_out <= x"600c0c05";
when 13 => instruction_out <= x"00004780";
when 14 => instruction_out <= x"400b0409";
when 15 => instruction_out <= x"00000780";
when 16 => instruction_out <= x"600a0609";
when 17 => instruction_out <= x"00008780";
when 18 => instruction_out <= x"30100409";
when 19 => instruction_out <= x"c4100780";
when 20 => instruction_out <= x"600a0405";
when 21 => instruction_out <= x"00008780";
when 22 => instruction_out <= x"a0004811";
when 23 => instruction_out <= x"04200780";
when 24 => instruction_out <= x"40090409";
when 25 => instruction_out <= x"00000780";
when 26 => instruction_out <= x"60080609";
when 27 => instruction_out <= x"00008780";
when 28 => instruction_out <= x"30100409";
when 29 => instruction_out <= x"c4100780";
when 30 => instruction_out <= x"60080421";
when 31 => instruction_out <= x"00008780";
when 32 => instruction_out <= x"1100ee04";
when 33 => instruction_out <= x"1100ec08";
when 34 => instruction_out <= x"a0004a1d";
when 35 => instruction_out <= x"04200780";
when 36 => instruction_out <= x"40050424";
when 37 => instruction_out <= x"40111c28";
when 38 => instruction_out <= x"60040625";
when 39 => instruction_out <= x"00024780";
when 40 => instruction_out <= x"60101e29";
when 41 => instruction_out <= x"00028780";
when 42 => instruction_out <= x"30101225";
when 43 => instruction_out <= x"c4100780";
when 44 => instruction_out <= x"30101429";
when 45 => instruction_out <= x"c4100780";
when 46 => instruction_out <= x"60040409";
when 47 => instruction_out <= x"00024780";
when 48 => instruction_out <= x"60101c05";
when 49 => instruction_out <= x"00028780";
when 50 => instruction_out <= x"307c05fd";
when 51 => instruction_out <= x"6c00c7c8";
when 52 => instruction_out <= x"10021003";
when 53 => instruction_out <= x"00000280";
when 54 => instruction_out <= x"1000f825";
when 55 => instruction_out <= x"0403c780";
when 56 => instruction_out <= x"30010409";
when 57 => instruction_out <= x"ec100780";
when 58 => instruction_out <= x"307c05fd";
when 59 => instruction_out <= x"6c0107c8";
when 60 => instruction_out <= x"20019225";
when 61 => instruction_out <= x"00000003";
when 62 => instruction_out <= x"1001c003";
when 63 => instruction_out <= x"00000280";
when 64 => instruction_out <= x"10022003";
when 65 => instruction_out <= x"00000780";
when 66 => instruction_out <= x"1000f825";
when 67 => instruction_out <= x"0403c780";
when 68 => instruction_out <= x"307c03fd";
when 69 => instruction_out <= x"6c00c7c8";
when 70 => instruction_out <= x"1002a003";
when 71 => instruction_out <= x"00000280";
when 72 => instruction_out <= x"1000f829";
when 73 => instruction_out <= x"0403c780";
when 74 => instruction_out <= x"30010205";
when 75 => instruction_out <= x"ec100780";
when 76 => instruction_out <= x"307c03fd";
when 77 => instruction_out <= x"6c0107c8";
when 78 => instruction_out <= x"20019429";
when 79 => instruction_out <= x"00000003";
when 80 => instruction_out <= x"10025003";
when 81 => instruction_out <= x"00000280";
when 82 => instruction_out <= x"1002b003";
when 83 => instruction_out <= x"00000780";
when 84 => instruction_out <= x"1000f829";
when 85 => instruction_out <= x"0403c780";
when 86 => instruction_out <= x"a0004e05";
when 87 => instruction_out <= x"04200780";
when 88 => instruction_out <= x"40021a09";
when 89 => instruction_out <= x"00000780";
when 90 => instruction_out <= x"60031809";
when 91 => instruction_out <= x"00008780";
when 92 => instruction_out <= x"30100409";
when 93 => instruction_out <= x"c4100780";
when 94 => instruction_out <= x"300a020d";
when 95 => instruction_out <= x"e0100780";
when 96 => instruction_out <= x"6002181d";
when 97 => instruction_out <= x"00008780";
when 98 => instruction_out <= x"a0004c09";
when 99 => instruction_out <= x"04200780";
when 100 => instruction_out <= x"a0000605";
when 101 => instruction_out <= x"04000780";
when 102 => instruction_out <= x"40021a20";
when 103 => instruction_out <= x"40041a2c";
when 104 => instruction_out <= x"400e0e31";
when 105 => instruction_out <= x"00000780";
when 106 => instruction_out <= x"60031821";
when 107 => instruction_out <= x"00020780";
when 108 => instruction_out <= x"6005182d";
when 109 => instruction_out <= x"0002c780";
when 110 => instruction_out <= x"600f0c31";
when 111 => instruction_out <= x"00030780";
when 112 => instruction_out <= x"30101021";
when 113 => instruction_out <= x"c4100780";
when 114 => instruction_out <= x"3010162d";
when 115 => instruction_out <= x"c4100780";
when 116 => instruction_out <= x"30101831";
when 117 => instruction_out <= x"c4100780";
when 118 => instruction_out <= x"60021805";
when 119 => instruction_out <= x"00020780";
when 120 => instruction_out <= x"60041809";
when 121 => instruction_out <= x"0002c780";
when 122 => instruction_out <= x"600e0c1d";
when 123 => instruction_out <= x"00030780";
when 124 => instruction_out <= x"d0800205";
when 125 => instruction_out <= x"00400780";
when 126 => instruction_out <= x"a0000221";
when 127 => instruction_out <= x"04000780";
when 128 => instruction_out <= x"40040e2d";
when 129 => instruction_out <= x"00000780";
when 130 => instruction_out <= x"400e1635";
when 131 => instruction_out <= x"00000780";
when 132 => instruction_out <= x"60050c31";
when 133 => instruction_out <= x"0002c780";
when 134 => instruction_out <= x"400d202d";
when 135 => instruction_out <= x"00000780";
when 136 => instruction_out <= x"600f143d";
when 137 => instruction_out <= x"00034780";
when 138 => instruction_out <= x"40070435";
when 139 => instruction_out <= x"00000780";
when 140 => instruction_out <= x"30101839";
when 141 => instruction_out <= x"c4100780";
when 142 => instruction_out <= x"600c2231";
when 143 => instruction_out <= x"0002c780";
when 144 => instruction_out <= x"30101e3d";
when 145 => instruction_out <= x"c4100780";
when 146 => instruction_out <= x"60060635";
when 147 => instruction_out <= x"00034780";
when 148 => instruction_out <= x"60040c2d";
when 149 => instruction_out <= x"00038780";
when 150 => instruction_out <= x"600e1409";
when 151 => instruction_out <= x"0003c780";
when 152 => instruction_out <= x"400b2c39";
when 153 => instruction_out <= x"00000780";
when 154 => instruction_out <= x"3010181d";
when 155 => instruction_out <= x"c4100780";
when 156 => instruction_out <= x"30101a31";
when 157 => instruction_out <= x"c4100780";
when 158 => instruction_out <= x"4009083d";
when 159 => instruction_out <= x"00000780";
when 160 => instruction_out <= x"600a2e35";
when 161 => instruction_out <= x"00038780";
when 162 => instruction_out <= x"600c2019";
when 163 => instruction_out <= x"0001c780";
when 164 => instruction_out <= x"6006040d";
when 165 => instruction_out <= x"00030780";
when 166 => instruction_out <= x"60080a21";
when 167 => instruction_out <= x"0003c780";
when 168 => instruction_out <= x"30101a1d";
when 169 => instruction_out <= x"c4100780";
when 170 => instruction_out <= x"204a9204";
when 171 => instruction_out <= x"20038c18";
when 172 => instruction_out <= x"30101021";
when 173 => instruction_out <= x"c4100780";
when 174 => instruction_out <= x"600a2c1d";
when 175 => instruction_out <= x"0001c780";
when 176 => instruction_out <= x"1001800d";
when 177 => instruction_out <= x"00000003";
when 178 => instruction_out <= x"a0000015";
when 179 => instruction_out <= x"04000780";
when 180 => instruction_out <= x"60080809";
when 181 => instruction_out <= x"00020780";
when 182 => instruction_out <= x"30010601";
when 183 => instruction_out <= x"c4000780";
when 184 => instruction_out <= x"20068a04";
when 185 => instruction_out <= x"20028e08";
when 186 => instruction_out <= x"3000cffd";
when 187 => instruction_out <= x"642047d8";
when 188 => instruction_out <= x"2000020d";
when 189 => instruction_out <= x"04008780";
when 190 => instruction_out <= x"307ccffd";
when 191 => instruction_out <= x"6c2107c8";
when 192 => instruction_out <= x"1009f003";
when 193 => instruction_out <= x"00001280";
when 194 => instruction_out <= x"1100ee04";
when 195 => instruction_out <= x"10008008";
when 196 => instruction_out <= x"10069003";
when 197 => instruction_out <= x"00000100";
when 198 => instruction_out <= x"1000f811";
when 199 => instruction_out <= x"0403c780";
when 200 => instruction_out <= x"30010205";
when 201 => instruction_out <= x"ec100780";
when 202 => instruction_out <= x"307c03fd";
when 203 => instruction_out <= x"6c0107d8";
when 204 => instruction_out <= x"20018811";
when 205 => instruction_out <= x"00000003";
when 206 => instruction_out <= x"10064003";
when 207 => instruction_out <= x"00001280";
when 208 => instruction_out <= x"1006a003";
when 209 => instruction_out <= x"00000780";
when 210 => instruction_out <= x"1000f811";
when 211 => instruction_out <= x"0403c780";
when 212 => instruction_out <= x"307c01fd";
when 213 => instruction_out <= x"6c00c7d8";
when 214 => instruction_out <= x"10072003";
when 215 => instruction_out <= x"00001280";
when 216 => instruction_out <= x"1000f805";
when 217 => instruction_out <= x"0403c780";
when 218 => instruction_out <= x"30010409";
when 219 => instruction_out <= x"ec100780";
when 220 => instruction_out <= x"307c05fd";
when 221 => instruction_out <= x"6c0107d8";
when 222 => instruction_out <= x"20018205";
when 223 => instruction_out <= x"00000003";
when 224 => instruction_out <= x"1006d003";
when 225 => instruction_out <= x"00001280";
when 226 => instruction_out <= x"10073003";
when 227 => instruction_out <= x"00000780";
when 228 => instruction_out <= x"1000f805";
when 229 => instruction_out <= x"0403c780";
when 230 => instruction_out <= x"20400805";
when 231 => instruction_out <= x"04004780";
when 232 => instruction_out <= x"10018009";
when 233 => instruction_out <= x"00000003";
when 234 => instruction_out <= x"30010409";
when 235 => instruction_out <= x"c4000780";
when 236 => instruction_out <= x"307c0405";
when 237 => instruction_out <= x"6c0107e0";
when 238 => instruction_out <= x"a00003fd";
when 239 => instruction_out <= x"0c0147d8";
when 240 => instruction_out <= x"10000405";
when 241 => instruction_out <= x"0403c780";
when 242 => instruction_out <= x"10080003";
when 243 => instruction_out <= x"00002100";
when 244 => instruction_out <= x"1000f811";
when 245 => instruction_out <= x"0403c780";
when 246 => instruction_out <= x"30010409";
when 247 => instruction_out <= x"ec100780";
when 248 => instruction_out <= x"307c05fd";
when 249 => instruction_out <= x"6c0107e8";
when 250 => instruction_out <= x"20018811";
when 251 => instruction_out <= x"00000003";
when 252 => instruction_out <= x"1007b003";
when 253 => instruction_out <= x"00002280";
when 254 => instruction_out <= x"10081003";
when 255 => instruction_out <= x"00000780";
when 256 => instruction_out <= x"1000f811";
when 257 => instruction_out <= x"0403c780";
when 258 => instruction_out <= x"203f8209";
when 259 => instruction_out <= x"0fffffff";
when 260 => instruction_out <= x"d0020615";
when 261 => instruction_out <= x"04000780";
when 262 => instruction_out <= x"400b0009";
when 263 => instruction_out <= x"00000780";
when 264 => instruction_out <= x"600a0219";
when 265 => instruction_out <= x"00008780";
when 266 => instruction_out <= x"203f8809";
when 267 => instruction_out <= x"0fffffff";
when 268 => instruction_out <= x"30100c11";
when 269 => instruction_out <= x"c4100780";
when 270 => instruction_out <= x"3002060d";
when 271 => instruction_out <= x"ec000780";
when 272 => instruction_out <= x"600a0011";
when 273 => instruction_out <= x"00010780";
when 274 => instruction_out <= x"1000ce01";
when 275 => instruction_out <= x"0423c780";
when 276 => instruction_out <= x"10091003";
when 277 => instruction_out <= x"00000100";
when 278 => instruction_out <= x"1000f809";
when 279 => instruction_out <= x"0403c780";
when 280 => instruction_out <= x"30010001";
when 281 => instruction_out <= x"ec100780";
when 282 => instruction_out <= x"307c01fd";
when 283 => instruction_out <= x"6c0107c8";
when 284 => instruction_out <= x"20018409";
when 285 => instruction_out <= x"00000003";
when 286 => instruction_out <= x"1008c003";
when 287 => instruction_out <= x"00000280";
when 288 => instruction_out <= x"10092003";
when 289 => instruction_out <= x"00000780";
when 290 => instruction_out <= x"1000f809";
when 291 => instruction_out <= x"0403c780";
when 292 => instruction_out <= x"10099003";
when 293 => instruction_out <= x"00001100";
when 294 => instruction_out <= x"1000f801";
when 295 => instruction_out <= x"0403c780";
when 296 => instruction_out <= x"30010205";
when 297 => instruction_out <= x"ec100780";
when 298 => instruction_out <= x"307c03fd";
when 299 => instruction_out <= x"6c0107c8";
when 300 => instruction_out <= x"20018001";
when 301 => instruction_out <= x"00000003";
when 302 => instruction_out <= x"10094003";
when 303 => instruction_out <= x"00000280";
when 304 => instruction_out <= x"1009a003";
when 305 => instruction_out <= x"00000780";
when 306 => instruction_out <= x"1000f801";
when 307 => instruction_out <= x"0403c780";
when 308 => instruction_out <= x"20400401";
when 309 => instruction_out <= x"04000780";
when 310 => instruction_out <= x"10018005";
when 311 => instruction_out <= x"00000003";
when 312 => instruction_out <= x"30000201";
when 313 => instruction_out <= x"c4000780";
when 314 => instruction_out <= x"10018015";
when 315 => instruction_out <= x"00000003";
when 316 => instruction_out <= x"100d8003";
when 317 => instruction_out <= x"00000780";
when 318 => instruction_out <= x"307c01fd";
when 319 => instruction_out <= x"6c00c7d8";
when 320 => instruction_out <= x"1000ce05";
when 321 => instruction_out <= x"0423c780";
when 322 => instruction_out <= x"100a8003";
when 323 => instruction_out <= x"00001280";
when 324 => instruction_out <= x"1000f809";
when 325 => instruction_out <= x"0403c780";
when 326 => instruction_out <= x"30010001";
when 327 => instruction_out <= x"ec100780";
when 328 => instruction_out <= x"307c01fd";
when 329 => instruction_out <= x"6c0107d8";
when 330 => instruction_out <= x"20018409";
when 331 => instruction_out <= x"00000003";
when 332 => instruction_out <= x"100a3003";
when 333 => instruction_out <= x"00001280";
when 334 => instruction_out <= x"100a9003";
when 335 => instruction_out <= x"00000780";
when 336 => instruction_out <= x"1000f809";
when 337 => instruction_out <= x"0403c780";
when 338 => instruction_out <= x"100b0003";
when 339 => instruction_out <= x"00000100";
when 340 => instruction_out <= x"1000f801";
when 341 => instruction_out <= x"0403c780";
when 342 => instruction_out <= x"30010205";
when 343 => instruction_out <= x"ec100780";
when 344 => instruction_out <= x"307c03fd";
when 345 => instruction_out <= x"6c0107c8";
when 346 => instruction_out <= x"20018001";
when 347 => instruction_out <= x"00000003";
when 348 => instruction_out <= x"100ab003";
when 349 => instruction_out <= x"00000280";
when 350 => instruction_out <= x"100b1003";
when 351 => instruction_out <= x"00000780";
when 352 => instruction_out <= x"1000f801";
when 353 => instruction_out <= x"0403c780";
when 354 => instruction_out <= x"20400401";
when 355 => instruction_out <= x"04000780";
when 356 => instruction_out <= x"10018005";
when 357 => instruction_out <= x"00000003";
when 358 => instruction_out <= x"30000205";
when 359 => instruction_out <= x"c4000780";
when 360 => instruction_out <= x"307c0201";
when 361 => instruction_out <= x"6c0107d0";
when 362 => instruction_out <= x"a00001fd";
when 363 => instruction_out <= x"0c0147c8";
when 364 => instruction_out <= x"10000201";
when 365 => instruction_out <= x"0403c780";
when 366 => instruction_out <= x"100be003";
when 367 => instruction_out <= x"00001100";
when 368 => instruction_out <= x"1000f809";
when 369 => instruction_out <= x"0403c780";
when 370 => instruction_out <= x"30010205";
when 371 => instruction_out <= x"ec100780";
when 372 => instruction_out <= x"307c03fd";
when 373 => instruction_out <= x"6c0107d8";
when 374 => instruction_out <= x"20018409";
when 375 => instruction_out <= x"00000003";
when 376 => instruction_out <= x"100b9003";
when 377 => instruction_out <= x"00001280";
when 378 => instruction_out <= x"100bf003";
when 379 => instruction_out <= x"00000780";
when 380 => instruction_out <= x"1000f809";
when 381 => instruction_out <= x"0403c780";
when 382 => instruction_out <= x"203f8405";
when 383 => instruction_out <= x"0fffffff";
when 384 => instruction_out <= x"307ccdfd";
when 385 => instruction_out <= x"6c20c7d8";
when 386 => instruction_out <= x"3001060d";
when 387 => instruction_out <= x"c4000780";
when 388 => instruction_out <= x"1000cc05";
when 389 => instruction_out <= x"0423c780";
when 390 => instruction_out <= x"100ca003";
when 391 => instruction_out <= x"00001280";
when 392 => instruction_out <= x"1000f809";
when 393 => instruction_out <= x"0403c780";
when 394 => instruction_out <= x"30010205";
when 395 => instruction_out <= x"ec100780";
when 396 => instruction_out <= x"307c03fd";
when 397 => instruction_out <= x"6c0107d8";
when 398 => instruction_out <= x"20018409";
when 399 => instruction_out <= x"00000003";
when 400 => instruction_out <= x"100c5003";
when 401 => instruction_out <= x"00001280";
when 402 => instruction_out <= x"100cb003";
when 403 => instruction_out <= x"00000780";
when 404 => instruction_out <= x"1000f809";
when 405 => instruction_out <= x"0403c780";
when 406 => instruction_out <= x"100d2003";
when 407 => instruction_out <= x"00000100";
when 408 => instruction_out <= x"1000f805";
when 409 => instruction_out <= x"0403c780";
when 410 => instruction_out <= x"30010001";
when 411 => instruction_out <= x"ec100780";
when 412 => instruction_out <= x"307c01fd";
when 413 => instruction_out <= x"6c0107c8";
when 414 => instruction_out <= x"20018205";
when 415 => instruction_out <= x"00000003";
when 416 => instruction_out <= x"100cd003";
when 417 => instruction_out <= x"00000280";
when 418 => instruction_out <= x"100d3003";
when 419 => instruction_out <= x"00000780";
when 420 => instruction_out <= x"1000f805";
when 421 => instruction_out <= x"0403c780";
when 422 => instruction_out <= x"20400401";
when 423 => instruction_out <= x"04004780";
when 424 => instruction_out <= x"10018005";
when 425 => instruction_out <= x"00000003";
when 426 => instruction_out <= x"30000215";
when 427 => instruction_out <= x"c4000780";
when 428 => instruction_out <= x"1000ce01";
when 429 => instruction_out <= x"0423c780";
when 430 => instruction_out <= x"1000f811";
when 431 => instruction_out <= x"0403c780";
when 432 => instruction_out <= x"307c0a05";
when 433 => instruction_out <= x"6c0107d0";
when 434 => instruction_out <= x"a00003fd";
when 435 => instruction_out <= x"0c0147c8";
when 436 => instruction_out <= x"10109003";
when 437 => instruction_out <= x"00001100";
when 438 => instruction_out <= x"307c01fd";
when 439 => instruction_out <= x"6c0107d8";
when 440 => instruction_out <= x"1000f821";
when 441 => instruction_out <= x"0403c780";
when 442 => instruction_out <= x"10106003";
when 443 => instruction_out <= x"00001100";
when 444 => instruction_out <= x"30040605";
when 445 => instruction_out <= x"c4100780";
when 446 => instruction_out <= x"30050609";
when 447 => instruction_out <= x"c4100780";
when 448 => instruction_out <= x"30010819";
when 449 => instruction_out <= x"c4100780";
when 450 => instruction_out <= x"20028208";
when 451 => instruction_out <= x"2006881c";
when 452 => instruction_out <= x"2000c809";
when 453 => instruction_out <= x"04208780";
when 454 => instruction_out <= x"30041019";
when 455 => instruction_out <= x"c4100780";
when 456 => instruction_out <= x"30051025";
when 457 => instruction_out <= x"c4100780";
when 458 => instruction_out <= x"20078408";
when 459 => instruction_out <= x"20018804";
when 460 => instruction_out <= x"20000c1d";
when 461 => instruction_out <= x"04024780";
when 462 => instruction_out <= x"30010029";
when 463 => instruction_out <= x"c4100780";
when 464 => instruction_out <= x"20068204";
when 465 => instruction_out <= x"20078424";
when 466 => instruction_out <= x"20001409";
when 467 => instruction_out <= x"04000780";
when 468 => instruction_out <= x"a0105003";
when 469 => instruction_out <= x"00000000";
when 470 => instruction_out <= x"21000229";
when 471 => instruction_out <= x"04408780";
when 472 => instruction_out <= x"2000122d";
when 473 => instruction_out <= x"04008780";
when 474 => instruction_out <= x"d00e1205";
when 475 => instruction_out <= x"80000780";
when 476 => instruction_out <= x"20019209";
when 477 => instruction_out <= x"00000003";
when 478 => instruction_out <= x"d00e0409";
when 479 => instruction_out <= x"80000780";
when 480 => instruction_out <= x"20029219";
when 481 => instruction_out <= x"00000003";
when 482 => instruction_out <= x"d00e0c1d";
when 483 => instruction_out <= x"80000780";
when 484 => instruction_out <= x"10058019";
when 485 => instruction_out <= x"00000967";
when 486 => instruction_out <= x"40041a31";
when 487 => instruction_out <= x"00000780";
when 488 => instruction_out <= x"30101831";
when 489 => instruction_out <= x"c4100780";
when 490 => instruction_out <= x"40048505";
when 491 => instruction_out <= x"000004cb";
when 492 => instruction_out <= x"60041809";
when 493 => instruction_out <= x"00030780";
when 494 => instruction_out <= x"30100205";
when 495 => instruction_out <= x"ec100780";
when 496 => instruction_out <= x"30100409";
when 497 => instruction_out <= x"ec100780";
when 498 => instruction_out <= x"401f9d19";
when 499 => instruction_out <= x"0000012f";
when 500 => instruction_out <= x"20000205";
when 501 => instruction_out <= x"04008780";
when 502 => instruction_out <= x"30100c09";
when 503 => instruction_out <= x"ec100780";
when 504 => instruction_out <= x"20000205";
when 505 => instruction_out <= x"04008780";
when 506 => instruction_out <= x"a0000405";
when 507 => instruction_out <= x"0c010780";
when 508 => instruction_out <= x"308103fd";
when 509 => instruction_out <= x"6c4107e8";
when 510 => instruction_out <= x"10000205";
when 511 => instruction_out <= x"2440e280";
when 512 => instruction_out <= x"20039225";
when 513 => instruction_out <= x"00000003";
when 514 => instruction_out <= x"d00e1405";
when 515 => instruction_out <= x"a0000780";
when 516 => instruction_out <= x"300b13fd";
when 517 => instruction_out <= x"640147e8";
when 518 => instruction_out <= x"20019429";
when 519 => instruction_out <= x"00000003";
when 520 => instruction_out <= x"100ed003";
when 521 => instruction_out <= x"00002280";
when 522 => instruction_out <= x"f0000001";
when 523 => instruction_out <= x"e0000002";
when 524 => instruction_out <= x"20019021";
when 525 => instruction_out <= x"00000003";
when 526 => instruction_out <= x"300511fd";
when 527 => instruction_out <= x"6c0147e8";
when 528 => instruction_out <= x"100dd003";
when 529 => instruction_out <= x"00002280";
when 530 => instruction_out <= x"30000003";
when 531 => instruction_out <= x"00000100";
when 532 => instruction_out <= x"307c01fd";
when 533 => instruction_out <= x"6c0107c8";
when 534 => instruction_out <= x"1000f819";
when 535 => instruction_out <= x"0403c780";
when 536 => instruction_out <= x"10160003";
when 537 => instruction_out <= x"00000100";
when 538 => instruction_out <= x"20018605";
when 539 => instruction_out <= x"00000003";
when 540 => instruction_out <= x"203f861d";
when 541 => instruction_out <= x"0fffffff";
when 542 => instruction_out <= x"213fec09";
when 543 => instruction_out <= x"0fffffff";
when 544 => instruction_out <= x"20018c04";
when 545 => instruction_out <= x"20078c1c";
when 546 => instruction_out <= x"300203fd";
when 547 => instruction_out <= x"6400c7d8";
when 548 => instruction_out <= x"307c0ffd";
when 549 => instruction_out <= x"6c0187e8";
when 550 => instruction_out <= x"a015f003";
when 551 => instruction_out <= x"00000000";
when 552 => instruction_out <= x"3004061d";
when 553 => instruction_out <= x"c4100780";
when 554 => instruction_out <= x"30040c21";
when 555 => instruction_out <= x"c4100780";
when 556 => instruction_out <= x"20018829";
when 557 => instruction_out <= x"00000003";
when 558 => instruction_out <= x"2104ea04";
when 559 => instruction_out <= x"20048e08";
when 560 => instruction_out <= x"213fee25";
when 561 => instruction_out <= x"0fffffff";
when 562 => instruction_out <= x"203f8831";
when 563 => instruction_out <= x"0fffffff";
when 564 => instruction_out <= x"20018e04";
when 565 => instruction_out <= x"20029008";
when 566 => instruction_out <= x"1000f83d";
when 567 => instruction_out <= x"0403c780";
when 568 => instruction_out <= x"2000942c";
when 569 => instruction_out <= x"20019034";
when 570 => instruction_out <= x"21000439";
when 571 => instruction_out <= x"04408780";
when 572 => instruction_out <= x"d00e1c05";
when 573 => instruction_out <= x"80000780";
when 574 => instruction_out <= x"403c8505";
when 575 => instruction_out <= x"0fffffff";
when 576 => instruction_out <= x"a0000405";
when 577 => instruction_out <= x"0c010780";
when 578 => instruction_out <= x"a012c003";
when 579 => instruction_out <= x"00000000";
when 580 => instruction_out <= x"300915fd";
when 581 => instruction_out <= x"640107f8";
when 582 => instruction_out <= x"1012c003";
when 583 => instruction_out <= x"00003280";
when 584 => instruction_out <= x"20049e08";
when 585 => instruction_out <= x"20079040";
when 586 => instruction_out <= x"20000409";
when 587 => instruction_out <= x"04040780";
when 588 => instruction_out <= x"21000409";
when 589 => instruction_out <= x"04408780";
when 590 => instruction_out <= x"20018409";
when 591 => instruction_out <= x"00000003";
when 592 => instruction_out <= x"d00e0409";
when 593 => instruction_out <= x"80000780";
when 594 => instruction_out <= x"a0000809";
when 595 => instruction_out <= x"04008780";
when 596 => instruction_out <= x"20000205";
when 597 => instruction_out <= x"04008780";
when 598 => instruction_out <= x"a0000405";
when 599 => instruction_out <= x"0c010780";
when 600 => instruction_out <= x"f0000001";
when 601 => instruction_out <= x"e0000002";
when 602 => instruction_out <= x"a0137003";
when 603 => instruction_out <= x"00000000";
when 604 => instruction_out <= x"10137003";
when 605 => instruction_out <= x"00001100";
when 606 => instruction_out <= x"20049e08";
when 607 => instruction_out <= x"20079040";
when 608 => instruction_out <= x"20000409";
when 609 => instruction_out <= x"04040780";
when 610 => instruction_out <= x"21000409";
when 611 => instruction_out <= x"04408780";
when 612 => instruction_out <= x"20108409";
when 613 => instruction_out <= x"00000003";
when 614 => instruction_out <= x"d00e0409";
when 615 => instruction_out <= x"80000780";
when 616 => instruction_out <= x"a0000809";
when 617 => instruction_out <= x"04008780";
when 618 => instruction_out <= x"20000205";
when 619 => instruction_out <= x"04008780";
when 620 => instruction_out <= x"a0000405";
when 621 => instruction_out <= x"0c010780";
when 622 => instruction_out <= x"f0000001";
when 623 => instruction_out <= x"e0000002";
when 624 => instruction_out <= x"a0143003";
when 625 => instruction_out <= x"00000000";
when 626 => instruction_out <= x"307c19fd";
when 627 => instruction_out <= x"6c0047f8";
when 628 => instruction_out <= x"10143003";
when 629 => instruction_out <= x"00003280";
when 630 => instruction_out <= x"20049e08";
when 631 => instruction_out <= x"20079040";
when 632 => instruction_out <= x"20000409";
when 633 => instruction_out <= x"04040780";
when 634 => instruction_out <= x"21000409";
when 635 => instruction_out <= x"04408780";
when 636 => instruction_out <= x"203f8409";
when 637 => instruction_out <= x"0fffffff";
when 638 => instruction_out <= x"d00e0409";
when 639 => instruction_out <= x"80000780";
when 640 => instruction_out <= x"a0000809";
when 641 => instruction_out <= x"04008780";
when 642 => instruction_out <= x"20000205";
when 643 => instruction_out <= x"04008780";
when 644 => instruction_out <= x"a0000405";
when 645 => instruction_out <= x"0c010780";
when 646 => instruction_out <= x"f0000001";
when 647 => instruction_out <= x"e0000002";
when 648 => instruction_out <= x"a014e003";
when 649 => instruction_out <= x"00000000";
when 650 => instruction_out <= x"1014e003";
when 651 => instruction_out <= x"00002100";
when 652 => instruction_out <= x"20049e08";
when 653 => instruction_out <= x"20079040";
when 654 => instruction_out <= x"20000409";
when 655 => instruction_out <= x"04040780";
when 656 => instruction_out <= x"21000409";
when 657 => instruction_out <= x"04408780";
when 658 => instruction_out <= x"20308409";
when 659 => instruction_out <= x"0fffffff";
when 660 => instruction_out <= x"d00e0409";
when 661 => instruction_out <= x"80000780";
when 662 => instruction_out <= x"a0000809";
when 663 => instruction_out <= x"04008780";
when 664 => instruction_out <= x"20000205";
when 665 => instruction_out <= x"04008780";
when 666 => instruction_out <= x"a0000405";
when 667 => instruction_out <= x"0c010780";
when 668 => instruction_out <= x"f0000001";
when 669 => instruction_out <= x"e0000002";
when 670 => instruction_out <= x"a0156003";
when 671 => instruction_out <= x"00000000";
when 672 => instruction_out <= x"307c03fd";
when 673 => instruction_out <= x"6c0187f8";
when 674 => instruction_out <= x"10154003";
when 675 => instruction_out <= x"00003280";
when 676 => instruction_out <= x"1000f805";
when 677 => instruction_out <= x"0403c780";
when 678 => instruction_out <= x"10156003";
when 679 => instruction_out <= x"00000780";
when 680 => instruction_out <= x"308103fd";
when 681 => instruction_out <= x"6c40c7f8";
when 682 => instruction_out <= x"10000205";
when 683 => instruction_out <= x"2440f500";
when 684 => instruction_out <= x"f0000001";
when 685 => instruction_out <= x"e0000002";
when 686 => instruction_out <= x"d00e1a05";
when 687 => instruction_out <= x"a0000780";
when 688 => instruction_out <= x"20019e3d";
when 689 => instruction_out <= x"00000003";
when 690 => instruction_out <= x"20019429";
when 691 => instruction_out <= x"00000003";
when 692 => instruction_out <= x"20019c39";
when 693 => instruction_out <= x"00000003";
when 694 => instruction_out <= x"20019831";
when 695 => instruction_out <= x"00000003";
when 696 => instruction_out <= x"20019a35";
when 697 => instruction_out <= x"00000003";
when 698 => instruction_out <= x"300b15fd";
when 699 => instruction_out <= x"6c0147f8";
when 700 => instruction_out <= x"1011e003";
when 701 => instruction_out <= x"00003280";
when 702 => instruction_out <= x"f0000001";
when 703 => instruction_out <= x"e0000002";
when 704 => instruction_out <= x"20018c19";
when 705 => instruction_out <= x"00000003";
when 706 => instruction_out <= x"30050dfd";
when 707 => instruction_out <= x"6c0147d8";
when 708 => instruction_out <= x"1010c003";
when 709 => instruction_out <= x"00001280";
when 710 => instruction_out <= x"f0000001";
when 711 => instruction_out <= x"e0000001";
when 712 => instruction_out <= x"30000003";
when 713 => instruction_out <= x"00000780";

			when others => null;
		end case;
	end process;

end arch;
