library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C0_reci is
	generic(
		word_bits	:natural:=26;
		bus_bits	:natural:=29;
		add_bits	:natural:=7
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C0_reci is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"11111111111111111111111110",
		"11111100000001111110111110",
		"11111000000111111000000110",
		"11110100010001100101100100",
		"11110000011111000001111010",
		"11101100110000000111101010",
		"11101001000100110001101000",
		"11100101011100111010110000",
		"11100001111000011110000100",
		"11011110010111010110110110",
		"11011010111001100000011100",
		"11010111011110110110010010",
		"11010100000111010100000100",
		"11010000110010110101100010",
		"11001101100001010110100000",
		"11001010010010110011000000",
		"11000111000111000111000100",
		"11000011111110001110111110",
		"11000000111000000110111110",
		"10111101110100101011100000",
		"10111010110011111001000100",
		"10110111110101101100001110",
		"10110100111010000001101100",
		"10110010000000110110001110",
		"10101111001010000110101110",
		"10101100010101110000000100",
		"10101001100011101111010110",
		"10100110110100000001101000",
		"10100100000110100100000100",
		"10100001011011010011111100",
		"10011110110010001110100100",
		"10011100001011010001010010",
		"10011001100110011001100100",
		"10010111000011100100111100",
		"10010100100010110000111110",
		"10010010000011111011010000",
		"10001111100111000001100010",
		"10001101001100000001100010",
		"10001010110010111001000010",
		"10001000011011100101111010",
		"10000110000110000110000100",
		"10000011110010010111011110",
		"10000001100000011000000100",
		"01111111010000000101111110",
		"01111101000001011111001110",
		"01111010110100100010000000",
		"01111000101001001100011110",
		"01110110011111011100111000",
		"01110100010111010001011100",
		"01110010010000101000011110",
		"01110000001011100000010110",
		"01101110000111110111011010",
		"01101100000101101100000100",
		"01101010000100111100110010",
		"01101000000101101000000100",
		"01100110000111101100011010",
		"01100100001011001000010100",
		"01100010001111111010011100",
		"01100000010110000001010110",
		"01011110011101011011101100",
		"01011100100110001000001010",
		"01011010110000000101011010",
		"01011000111011010010001010",
		"01010111000111101101001110",
		"01010101010101010101010100",
		"01010011100100001001010000",
		"01010001110100000111111010",
		"01010000000101010000000100",
		"01001110010111100000101000",
		"01001100101010111000100000",
		"01001010111111010110100110",
		"01001001010100111001111000",
		"01000111101011100001010000",
		"01000110000011001011110000",
		"01000100011011111000011000",
		"01000010110101100110001000",
		"01000001010000010100000100",
		"00111111101100000001001110",
		"00111110001000101100101110",
		"00111100100110010101101000",
		"00111011000100111011000100",
		"00111001100100011100001010",
		"00111000000100111000000100",
		"00110110100110001101111100",
		"00110101001000011100111110",
		"00110011101011100100010110",
		"00110010001111100011010010",
		"00110000110100011001000000",
		"00101111011010000100101110",
		"00101110000000100101101110",
		"00101100100111111011010010",
		"00101011010000000100101010",
		"00101001111001000001001010",
		"00101000100010110000000100",
		"00100111001101010000101100",
		"00100101111000100010011010",
		"00100100100100100100100100",
		"00100011010001010110011100",
		"00100001111110110111100000",
		"00100000101101000111000010",
		"00011111011100000100011110",
		"00011110001011101111001110",
		"00011100111100000110101010",
		"00011011101101001010001110",
		"00011010011110111001011000",
		"00011001010001010011011110",
		"00011000000100011000000100",
		"00010110111000000110100010",
		"00010101101100011110010110",
		"00010100100001011111000010",
		"00010011010111001000000100",
		"00010010001101011000111000",
		"00010001000100010001000100",
		"00001111111011110000000100",
		"00001110110011110101011010",
		"00001101101100100000101010",
		"00001100100101110001010010",
		"00001011011111100110111010",
		"00001010011010000001000010",
		"00001001010100111111001110",
		"00001000010000100001000000",
		"00000111001100100110000010",
		"00000110001001001101110100",
		"00000101000110010111111100",
		"00000100000100000100000010",
		"00000011000010010001101100",
		"00000010000001000000100000",
		"00000001000000010000000010"
	);
begin
	data <= "001"&rom(to_integer(unsigned(addr)));
end architecture;