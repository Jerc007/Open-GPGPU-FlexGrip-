library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LUT_C1_sqrt_2_4 is
	generic(
		word_bits	:natural:=16;
		bus_bits	:natural:=20;
		add_bits	:natural:=6
	);
	port(
		addr		:in std_logic_vector(add_bits-1 downto 0);
		data		:out std_logic_vector(bus_bits-1 downto 0)
	);
end entity;

architecture behav of LUT_C1_sqrt_2_4 is
	type storage is array (0 to 2**add_bits-1) of std_logic_vector(word_bits-1 downto 0);
	constant rom:storage:=(
		"1101010000010000",
		"1100111001111000",
		"1100100100000000",
		"1100001110101000",
		"1011111001110000",
		"1011100101010000",
		"1011010001010000",
		"1010111101110000",
		"1010101010101000",
		"1010010111110000",
		"1010000101011000",
		"1001110011011000",
		"1001100001110000",
		"1001010000011000",
		"1000111111100000",
		"1000101110110000",
		"1000011110100000",
		"1000001110011000",
		"0111111110101000",
		"0111101111010000",
		"0111100000000000",
		"0111010001001000",
		"0111000010100000",
		"0110110100000000",
		"0110100101111000",
		"0110011000000000",
		"0110001010010000",
		"0101111100111000",
		"0101101111101000",
		"0101100010101000",
		"0101010101110000",
		"0101001001001000",
		"0100111100110000",
		"0100110000100000",
		"0100100100100000",
		"0100011000101000",
		"0100001101000000",
		"0100000001100000",
		"0011110110001000",
		"0011101011000000",
		"0011100000000000",
		"0011010101001000",
		"0011001010100000",
		"0010111111111000",
		"0010110101100000",
		"0010101011010000",
		"0010100001001000",
		"0010010111001000",
		"0010001101011000",
		"0010000011101000",
		"0001111010000000",
		"0001110000101000",
		"0001100111010000",
		"0001011110000000",
		"0001010101000000",
		"0001001100000000",
		"0001000011001000",
		"0000111010011000",
		"0000110001101000",
		"0000101001001000",
		"0000100000110000",
		"0000011000011000",
		"0000010000001000",
		"0000001000000000"
	);
begin
	data <= "0010"&rom(to_integer(unsigned(addr)));
end architecture;