
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity TP_instructions is
	port(
		instruction_pointer_in : in  integer;
		num_instructions_out   : out integer;
		instruction_out        : out std_logic_vector(31 downto 0)
	);
end TP_instructions;

architecture arch of TP_instructions is
	constant TP_INSTRUCTIONS : integer := 786;

begin
	num_instructions_out <= TP_INSTRUCTIONS;

	process(instruction_pointer_in)
	begin
		case instruction_pointer_in is
			                when 0 => instruction_out <= x"10008028";   -- MOV32 R10, R0;
                when 1 => instruction_out <= x"10018031";   -- MVI R12, 0x1;
                when 2 => instruction_out <= x"00000003";
                when 3 => instruction_out <= x"300c1831";   -- SHL R12, R12, 0xc;
                when 4 => instruction_out <= x"c4100780";
                when 5 => instruction_out <= x"20009830";   -- IADD32 R12, R12, R0;
                when 6 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 7 => instruction_out <= x"80c00780";
                when 8 => instruction_out <= x"10008035";   -- MVI R13, 0x0;
                when 9 => instruction_out <= x"00000003";
                when 10 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 11 => instruction_out <= x"a0c00780";
                when 12 => instruction_out <= x"1001802d";   -- MVI R11, 0x1;
                when 13 => instruction_out <= x"00000003";
                when 14 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 15 => instruction_out <= x"040087c0";
                when 16 => instruction_out <= x"a0011003";   -- SSY 0x88;
                when 17 => instruction_out <= x"00000780";
                when 18 => instruction_out <= x"1000c003";   -- BRA (C48.EQU), 0x60;
                when 19 => instruction_out <= x"00000500";
                when 20 => instruction_out <= x"f0000001";   -- NOP;
                when 21 => instruction_out <= x"e0000000";
                when 22 => instruction_out <= x"10010003";   -- BRA 0x80;
                when 23 => instruction_out <= x"00000780";
                when 24 => instruction_out <= x"f0000001";   -- NOP;
                when 25 => instruction_out <= x"e0000000";
                when 26 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 27 => instruction_out <= x"80c00780";
                when 28 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 29 => instruction_out <= x"00000003";
                when 30 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 31 => instruction_out <= x"a0c00780";
                when 32 => instruction_out <= x"f0000001";   -- NOP;
                when 33 => instruction_out <= x"e0000000";
                when 34 => instruction_out <= x"f0000001";   -- NOP.S;
                when 35 => instruction_out <= x"e0000002";
                when 36 => instruction_out <= x"1002802d";   -- MVI R11, 0x2;
                when 37 => instruction_out <= x"00000003";
                when 38 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 39 => instruction_out <= x"040087c0";
                when 40 => instruction_out <= x"a001d003";   -- SSY 0xe8;
                when 41 => instruction_out <= x"00000780";
                when 42 => instruction_out <= x"10018003";   -- BRA (C48.EQU), 0xc0;
                when 43 => instruction_out <= x"00000500";
                when 44 => instruction_out <= x"f0000001";   -- NOP;
                when 45 => instruction_out <= x"e0000000";
                when 46 => instruction_out <= x"1001c003";   -- BRA 0xe0;
                when 47 => instruction_out <= x"00000780";
                when 48 => instruction_out <= x"f0000001";   -- NOP;
                when 49 => instruction_out <= x"e0000000";
                when 50 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 51 => instruction_out <= x"80c00780";
                when 52 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 53 => instruction_out <= x"00000003";
                when 54 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 55 => instruction_out <= x"a0c00780";
                when 56 => instruction_out <= x"f0000001";   -- NOP;
                when 57 => instruction_out <= x"e0000000";
                when 58 => instruction_out <= x"f0000001";   -- NOP.S;
                when 59 => instruction_out <= x"e0000002";
                when 60 => instruction_out <= x"1003802d";   -- MVI R11, 0x3;
                when 61 => instruction_out <= x"00000003";
                when 62 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 63 => instruction_out <= x"040087c0";
                when 64 => instruction_out <= x"a0029003";   -- SSY 0x148;
                when 65 => instruction_out <= x"00000780";
                when 66 => instruction_out <= x"10024003";   -- BRA (C48.EQU), 0x120;
                when 67 => instruction_out <= x"00000500";
                when 68 => instruction_out <= x"f0000001";   -- NOP;
                when 69 => instruction_out <= x"e0000000";
                when 70 => instruction_out <= x"10028003";   -- BRA 0x140;
                when 71 => instruction_out <= x"00000780";
                when 72 => instruction_out <= x"f0000001";   -- NOP;
                when 73 => instruction_out <= x"e0000000";
                when 74 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 75 => instruction_out <= x"80c00780";
                when 76 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 77 => instruction_out <= x"00000003";
                when 78 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 79 => instruction_out <= x"a0c00780";
                when 80 => instruction_out <= x"f0000001";   -- NOP;
                when 81 => instruction_out <= x"e0000000";
                when 82 => instruction_out <= x"f0000001";   -- NOP.S;
                when 83 => instruction_out <= x"e0000002";
                when 84 => instruction_out <= x"1004802d";   -- MVI R11, 0x4;
                when 85 => instruction_out <= x"00000003";
                when 86 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 87 => instruction_out <= x"040087c0";
                when 88 => instruction_out <= x"a0035003";   -- SSY 0x1a8;
                when 89 => instruction_out <= x"00000780";
                when 90 => instruction_out <= x"10030003";   -- BRA (C48.EQU), 0x180;
                when 91 => instruction_out <= x"00000500";
                when 92 => instruction_out <= x"f0000001";   -- NOP;
                when 93 => instruction_out <= x"e0000000";
                when 94 => instruction_out <= x"10034003";   -- BRA 0x1a0;
                when 95 => instruction_out <= x"00000780";
                when 96 => instruction_out <= x"f0000001";   -- NOP;
                when 97 => instruction_out <= x"e0000000";
                when 98 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 99 => instruction_out <= x"80c00780";
                when 100 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 101 => instruction_out <= x"00000003";
                when 102 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 103 => instruction_out <= x"a0c00780";
                when 104 => instruction_out <= x"f0000001";   -- NOP;
                when 105 => instruction_out <= x"e0000000";
                when 106 => instruction_out <= x"f0000001";   -- NOP.S;
                when 107 => instruction_out <= x"e0000002";
                when 108 => instruction_out <= x"1005802d";   -- MVI R11, 0x5;
                when 109 => instruction_out <= x"00000003";
                when 110 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 111 => instruction_out <= x"040087c0";
                when 112 => instruction_out <= x"a0041003";   -- SSY 0x208;
                when 113 => instruction_out <= x"00000780";
                when 114 => instruction_out <= x"1003c003";   -- BRA (C48.EQU), 0x1e0;
                when 115 => instruction_out <= x"00000500";
                when 116 => instruction_out <= x"f0000001";   -- NOP;
                when 117 => instruction_out <= x"e0000000";
                when 118 => instruction_out <= x"10040003";   -- BRA 0x200;
                when 119 => instruction_out <= x"00000780";
                when 120 => instruction_out <= x"f0000001";   -- NOP;
                when 121 => instruction_out <= x"e0000000";
                when 122 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 123 => instruction_out <= x"80c00780";
                when 124 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 125 => instruction_out <= x"00000003";
                when 126 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 127 => instruction_out <= x"a0c00780";
                when 128 => instruction_out <= x"f0000001";   -- NOP;
                when 129 => instruction_out <= x"e0000000";
                when 130 => instruction_out <= x"f0000001";   -- NOP.S;
                when 131 => instruction_out <= x"e0000002";
                when 132 => instruction_out <= x"1006802d";   -- MVI R11, 0x6;
                when 133 => instruction_out <= x"00000003";
                when 134 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 135 => instruction_out <= x"040087c0";
                when 136 => instruction_out <= x"a004d003";   -- SSY 0x268;
                when 137 => instruction_out <= x"00000780";
                when 138 => instruction_out <= x"10048003";   -- BRA (C48.EQU), 0x240;
                when 139 => instruction_out <= x"00000500";
                when 140 => instruction_out <= x"f0000001";   -- NOP;
                when 141 => instruction_out <= x"e0000000";
                when 142 => instruction_out <= x"1004c003";   -- BRA 0x260;
                when 143 => instruction_out <= x"00000780";
                when 144 => instruction_out <= x"f0000001";   -- NOP;
                when 145 => instruction_out <= x"e0000000";
                when 146 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 147 => instruction_out <= x"80c00780";
                when 148 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 149 => instruction_out <= x"00000003";
                when 150 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 151 => instruction_out <= x"a0c00780";
                when 152 => instruction_out <= x"f0000001";   -- NOP;
                when 153 => instruction_out <= x"e0000000";
                when 154 => instruction_out <= x"f0000001";   -- NOP.S;
                when 155 => instruction_out <= x"e0000002";
                when 156 => instruction_out <= x"1007802d";   -- MVI R11, 0x7;
                when 157 => instruction_out <= x"00000003";
                when 158 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 159 => instruction_out <= x"040087c0";
                when 160 => instruction_out <= x"a0059003";   -- SSY 0x2c8;
                when 161 => instruction_out <= x"00000780";
                when 162 => instruction_out <= x"10054003";   -- BRA (C48.EQU), 0x2a0;
                when 163 => instruction_out <= x"00000500";
                when 164 => instruction_out <= x"f0000001";   -- NOP;
                when 165 => instruction_out <= x"e0000000";
                when 166 => instruction_out <= x"10058003";   -- BRA 0x2c0;
                when 167 => instruction_out <= x"00000780";
                when 168 => instruction_out <= x"f0000001";   -- NOP;
                when 169 => instruction_out <= x"e0000000";
                when 170 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 171 => instruction_out <= x"80c00780";
                when 172 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 173 => instruction_out <= x"00000003";
                when 174 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 175 => instruction_out <= x"a0c00780";
                when 176 => instruction_out <= x"f0000001";   -- NOP;
                when 177 => instruction_out <= x"e0000000";
                when 178 => instruction_out <= x"f0000001";   -- NOP.S;
                when 179 => instruction_out <= x"e0000002";
                when 180 => instruction_out <= x"1008802d";   -- MVI R11, 0x8;
                when 181 => instruction_out <= x"00000003";
                when 182 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 183 => instruction_out <= x"040087c0";
                when 184 => instruction_out <= x"a0065003";   -- SSY 0x328;
                when 185 => instruction_out <= x"00000780";
                when 186 => instruction_out <= x"10060003";   -- BRA (C48.EQU), 0x300;
                when 187 => instruction_out <= x"00000500";
                when 188 => instruction_out <= x"f0000001";   -- NOP;
                when 189 => instruction_out <= x"e0000000";
                when 190 => instruction_out <= x"10064003";   -- BRA 0x320;
                when 191 => instruction_out <= x"00000780";
                when 192 => instruction_out <= x"f0000001";   -- NOP;
                when 193 => instruction_out <= x"e0000000";
                when 194 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 195 => instruction_out <= x"80c00780";
                when 196 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 197 => instruction_out <= x"00000003";
                when 198 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 199 => instruction_out <= x"a0c00780";
                when 200 => instruction_out <= x"f0000001";   -- NOP;
                when 201 => instruction_out <= x"e0000000";
                when 202 => instruction_out <= x"f0000001";   -- NOP.S;
                when 203 => instruction_out <= x"e0000002";
                when 204 => instruction_out <= x"1009802d";   -- MVI R11, 0x9;
                when 205 => instruction_out <= x"00000003";
                when 206 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 207 => instruction_out <= x"040087c0";
                when 208 => instruction_out <= x"a0071003";   -- SSY 0x388;
                when 209 => instruction_out <= x"00000780";
                when 210 => instruction_out <= x"1006c003";   -- BRA (C48.EQU), 0x360;
                when 211 => instruction_out <= x"00000500";
                when 212 => instruction_out <= x"f0000001";   -- NOP;
                when 213 => instruction_out <= x"e0000000";
                when 214 => instruction_out <= x"10070003";   -- BRA 0x380;
                when 215 => instruction_out <= x"00000780";
                when 216 => instruction_out <= x"f0000001";   -- NOP;
                when 217 => instruction_out <= x"e0000000";
                when 218 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 219 => instruction_out <= x"80c00780";
                when 220 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 221 => instruction_out <= x"00000003";
                when 222 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 223 => instruction_out <= x"a0c00780";
                when 224 => instruction_out <= x"f0000001";   -- NOP;
                when 225 => instruction_out <= x"e0000000";
                when 226 => instruction_out <= x"f0000001";   -- NOP.S;
                when 227 => instruction_out <= x"e0000002";
                when 228 => instruction_out <= x"1009802d";   -- MVI R11, 0x9;
                when 229 => instruction_out <= x"00000003";
                when 230 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 231 => instruction_out <= x"040087c0";
                when 232 => instruction_out <= x"a007d003";   -- SSY 0x3e8;
                when 233 => instruction_out <= x"00000780";
                when 234 => instruction_out <= x"10078003";   -- BRA (C48.EQU), 0x3c0;
                when 235 => instruction_out <= x"00000500";
                when 236 => instruction_out <= x"f0000001";   -- NOP;
                when 237 => instruction_out <= x"e0000000";
                when 238 => instruction_out <= x"1007c003";   -- BRA 0x3e0;
                when 239 => instruction_out <= x"00000780";
                when 240 => instruction_out <= x"f0000001";   -- NOP;
                when 241 => instruction_out <= x"e0000000";
                when 242 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 243 => instruction_out <= x"80c00780";
                when 244 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 245 => instruction_out <= x"00000003";
                when 246 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 247 => instruction_out <= x"a0c00780";
                when 248 => instruction_out <= x"f0000001";   -- NOP;
                when 249 => instruction_out <= x"e0000000";
                when 250 => instruction_out <= x"f0000001";   -- NOP.S;
                when 251 => instruction_out <= x"e0000002";
                when 252 => instruction_out <= x"100a802d";   -- MVI R11, 0xa;
                when 253 => instruction_out <= x"00000003";
                when 254 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 255 => instruction_out <= x"040087c0";
                when 256 => instruction_out <= x"a0089003";   -- SSY 0x448;
                when 257 => instruction_out <= x"00000780";
                when 258 => instruction_out <= x"10084003";   -- BRA (C48.EQU), 0x420;
                when 259 => instruction_out <= x"00000500";
                when 260 => instruction_out <= x"f0000001";   -- NOP;
                when 261 => instruction_out <= x"e0000000";
                when 262 => instruction_out <= x"10088003";   -- BRA 0x440;
                when 263 => instruction_out <= x"00000780";
                when 264 => instruction_out <= x"f0000001";   -- NOP;
                when 265 => instruction_out <= x"e0000000";
                when 266 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 267 => instruction_out <= x"80c00780";
                when 268 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 269 => instruction_out <= x"00000003";
                when 270 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 271 => instruction_out <= x"a0c00780";
                when 272 => instruction_out <= x"f0000001";   -- NOP;
                when 273 => instruction_out <= x"e0000000";
                when 274 => instruction_out <= x"f0000001";   -- NOP.S;
                when 275 => instruction_out <= x"e0000002";
                when 276 => instruction_out <= x"100b802d";   -- MVI R11, 0xb;
                when 277 => instruction_out <= x"00000003";
                when 278 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 279 => instruction_out <= x"040087c0";
                when 280 => instruction_out <= x"a0095003";   -- SSY 0x4a8;
                when 281 => instruction_out <= x"00000780";
                when 282 => instruction_out <= x"10090003";   -- BRA (C48.EQU), 0x480;
                when 283 => instruction_out <= x"00000500";
                when 284 => instruction_out <= x"f0000001";   -- NOP;
                when 285 => instruction_out <= x"e0000000";
                when 286 => instruction_out <= x"10094003";   -- BRA 0x4a0;
                when 287 => instruction_out <= x"00000780";
                when 288 => instruction_out <= x"f0000001";   -- NOP;
                when 289 => instruction_out <= x"e0000000";
                when 290 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 291 => instruction_out <= x"80c00780";
                when 292 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 293 => instruction_out <= x"00000003";
                when 294 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 295 => instruction_out <= x"a0c00780";
                when 296 => instruction_out <= x"f0000001";   -- NOP;
                when 297 => instruction_out <= x"e0000000";
                when 298 => instruction_out <= x"f0000001";   -- NOP.S;
                when 299 => instruction_out <= x"e0000002";
                when 300 => instruction_out <= x"100c802d";   -- MVI R11, 0xc;
                when 301 => instruction_out <= x"00000003";
                when 302 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 303 => instruction_out <= x"040087c0";
                when 304 => instruction_out <= x"a00a1003";   -- SSY 0x508;
                when 305 => instruction_out <= x"00000780";
                when 306 => instruction_out <= x"1009c003";   -- BRA (C48.EQU), 0x4e0;
                when 307 => instruction_out <= x"00000500";
                when 308 => instruction_out <= x"f0000001";   -- NOP;
                when 309 => instruction_out <= x"e0000000";
                when 310 => instruction_out <= x"100a0003";   -- BRA 0x500;
                when 311 => instruction_out <= x"00000780";
                when 312 => instruction_out <= x"f0000001";   -- NOP;
                when 313 => instruction_out <= x"e0000000";
                when 314 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 315 => instruction_out <= x"80c00780";
                when 316 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 317 => instruction_out <= x"00000003";
                when 318 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 319 => instruction_out <= x"a0c00780";
                when 320 => instruction_out <= x"f0000001";   -- NOP;
                when 321 => instruction_out <= x"e0000000";
                when 322 => instruction_out <= x"f0000001";   -- NOP.S;
                when 323 => instruction_out <= x"e0000002";
                when 324 => instruction_out <= x"100d802d";   -- MVI R11, 0xd;
                when 325 => instruction_out <= x"00000003";
                when 326 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 327 => instruction_out <= x"040087c0";
                when 328 => instruction_out <= x"a00ad003";   -- SSY 0x568;
                when 329 => instruction_out <= x"00000780";
                when 330 => instruction_out <= x"100a8003";   -- BRA (C48.EQU), 0x540;
                when 331 => instruction_out <= x"00000500";
                when 332 => instruction_out <= x"f0000001";   -- NOP;
                when 333 => instruction_out <= x"e0000000";
                when 334 => instruction_out <= x"100ac003";   -- BRA 0x560;
                when 335 => instruction_out <= x"00000780";
                when 336 => instruction_out <= x"f0000001";   -- NOP;
                when 337 => instruction_out <= x"e0000000";
                when 338 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 339 => instruction_out <= x"80c00780";
                when 340 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 341 => instruction_out <= x"00000003";
                when 342 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 343 => instruction_out <= x"a0c00780";
                when 344 => instruction_out <= x"f0000001";   -- NOP;
                when 345 => instruction_out <= x"e0000000";
                when 346 => instruction_out <= x"f0000001";   -- NOP.S;
                when 347 => instruction_out <= x"e0000002";
                when 348 => instruction_out <= x"100e802d";   -- MVI R11, 0xe;
                when 349 => instruction_out <= x"00000003";
                when 350 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 351 => instruction_out <= x"040087c0";
                when 352 => instruction_out <= x"a00b9003";   -- SSY 0x5c8;
                when 353 => instruction_out <= x"00000780";
                when 354 => instruction_out <= x"100b4003";   -- BRA (C48.EQU), 0x5a0;
                when 355 => instruction_out <= x"00000500";
                when 356 => instruction_out <= x"f0000001";   -- NOP;
                when 357 => instruction_out <= x"e0000000";
                when 358 => instruction_out <= x"100b8003";   -- BRA 0x5c0;
                when 359 => instruction_out <= x"00000780";
                when 360 => instruction_out <= x"f0000001";   -- NOP;
                when 361 => instruction_out <= x"e0000000";
                when 362 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 363 => instruction_out <= x"80c00780";
                when 364 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 365 => instruction_out <= x"00000003";
                when 366 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 367 => instruction_out <= x"a0c00780";
                when 368 => instruction_out <= x"f0000001";   -- NOP;
                when 369 => instruction_out <= x"e0000000";
                when 370 => instruction_out <= x"f0000001";   -- NOP.S;
                when 371 => instruction_out <= x"e0000002";
                when 372 => instruction_out <= x"100f802d";   -- MVI R11, 0xf;
                when 373 => instruction_out <= x"00000003";
                when 374 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 375 => instruction_out <= x"040087c0";
                when 376 => instruction_out <= x"a00c5003";   -- SSY 0x628;
                when 377 => instruction_out <= x"00000780";
                when 378 => instruction_out <= x"100c0003";   -- BRA (C48.EQU), 0x600;
                when 379 => instruction_out <= x"00000500";
                when 380 => instruction_out <= x"f0000001";   -- NOP;
                when 381 => instruction_out <= x"e0000000";
                when 382 => instruction_out <= x"100c4003";   -- BRA 0x620;
                when 383 => instruction_out <= x"00000780";
                when 384 => instruction_out <= x"f0000001";   -- NOP;
                when 385 => instruction_out <= x"e0000000";
                when 386 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 387 => instruction_out <= x"80c00780";
                when 388 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 389 => instruction_out <= x"00000003";
                when 390 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 391 => instruction_out <= x"a0c00780";
                when 392 => instruction_out <= x"f0000001";   -- NOP;
                when 393 => instruction_out <= x"e0000000";
                when 394 => instruction_out <= x"f0000001";   -- NOP.S;
                when 395 => instruction_out <= x"e0000002";
                when 396 => instruction_out <= x"1010802d";   -- MVI R11, 0x10;
                when 397 => instruction_out <= x"00000003";
                when 398 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 399 => instruction_out <= x"040087c0";
                when 400 => instruction_out <= x"a00d1003";   -- SSY 0x688;
                when 401 => instruction_out <= x"00000780";
                when 402 => instruction_out <= x"100cc003";   -- BRA (C48.EQU), 0x660;
                when 403 => instruction_out <= x"00000500";
                when 404 => instruction_out <= x"f0000001";   -- NOP;
                when 405 => instruction_out <= x"e0000000";
                when 406 => instruction_out <= x"100d0003";   -- BRA 0x680;
                when 407 => instruction_out <= x"00000780";
                when 408 => instruction_out <= x"f0000001";   -- NOP;
                when 409 => instruction_out <= x"e0000000";
                when 410 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 411 => instruction_out <= x"80c00780";
                when 412 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 413 => instruction_out <= x"00000003";
                when 414 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 415 => instruction_out <= x"a0c00780";
                when 416 => instruction_out <= x"f0000001";   -- NOP;
                when 417 => instruction_out <= x"e0000000";
                when 418 => instruction_out <= x"f0000001";   -- NOP.S;
                when 419 => instruction_out <= x"e0000002";
                when 420 => instruction_out <= x"1011802d";   -- MVI R11, 0x11;
                when 421 => instruction_out <= x"00000003";
                when 422 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 423 => instruction_out <= x"040087c0";
                when 424 => instruction_out <= x"a00dd003";   -- SSY 0x6e8;
                when 425 => instruction_out <= x"00000780";
                when 426 => instruction_out <= x"100d8003";   -- BRA (C48.EQU), 0x6c0;
                when 427 => instruction_out <= x"00000500";
                when 428 => instruction_out <= x"f0000001";   -- NOP;
                when 429 => instruction_out <= x"e0000000";
                when 430 => instruction_out <= x"100dc003";   -- BRA 0x6e0;
                when 431 => instruction_out <= x"00000780";
                when 432 => instruction_out <= x"f0000001";   -- NOP;
                when 433 => instruction_out <= x"e0000000";
                when 434 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 435 => instruction_out <= x"80c00780";
                when 436 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 437 => instruction_out <= x"00000003";
                when 438 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 439 => instruction_out <= x"a0c00780";
                when 440 => instruction_out <= x"f0000001";   -- NOP;
                when 441 => instruction_out <= x"e0000000";
                when 442 => instruction_out <= x"f0000001";   -- NOP.S;
                when 443 => instruction_out <= x"e0000002";
                when 444 => instruction_out <= x"1012802d";   -- MVI R11, 0x12;
                when 445 => instruction_out <= x"00000003";
                when 446 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 447 => instruction_out <= x"040087c0";
                when 448 => instruction_out <= x"a00e9003";   -- SSY 0x748;
                when 449 => instruction_out <= x"00000780";
                when 450 => instruction_out <= x"100e4003";   -- BRA (C48.EQU), 0x720;
                when 451 => instruction_out <= x"00000500";
                when 452 => instruction_out <= x"f0000001";   -- NOP;
                when 453 => instruction_out <= x"e0000000";
                when 454 => instruction_out <= x"100e8003";   -- BRA 0x740;
                when 455 => instruction_out <= x"00000780";
                when 456 => instruction_out <= x"f0000001";   -- NOP;
                when 457 => instruction_out <= x"e0000000";
                when 458 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 459 => instruction_out <= x"80c00780";
                when 460 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 461 => instruction_out <= x"00000003";
                when 462 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 463 => instruction_out <= x"a0c00780";
                when 464 => instruction_out <= x"f0000001";   -- NOP;
                when 465 => instruction_out <= x"e0000000";
                when 466 => instruction_out <= x"f0000001";   -- NOP.S;
                when 467 => instruction_out <= x"e0000002";
                when 468 => instruction_out <= x"1013802d";   -- MVI R11, 0x13;
                when 469 => instruction_out <= x"00000003";
                when 470 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 471 => instruction_out <= x"040087c0";
                when 472 => instruction_out <= x"a00f5003";   -- SSY 0x7a8;
                when 473 => instruction_out <= x"00000780";
                when 474 => instruction_out <= x"100f0003";   -- BRA (C48.EQU), 0x780;
                when 475 => instruction_out <= x"00000500";
                when 476 => instruction_out <= x"f0000001";   -- NOP;
                when 477 => instruction_out <= x"e0000000";
                when 478 => instruction_out <= x"100f4003";   -- BRA 0x7a0;
                when 479 => instruction_out <= x"00000780";
                when 480 => instruction_out <= x"f0000001";   -- NOP;
                when 481 => instruction_out <= x"e0000000";
                when 482 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 483 => instruction_out <= x"80c00780";
                when 484 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 485 => instruction_out <= x"00000003";
                when 486 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 487 => instruction_out <= x"a0c00780";
                when 488 => instruction_out <= x"f0000001";   -- NOP;
                when 489 => instruction_out <= x"e0000000";
                when 490 => instruction_out <= x"f0000001";   -- NOP.S;
                when 491 => instruction_out <= x"e0000002";
                when 492 => instruction_out <= x"1014802d";   -- MVI R11, 0x14;
                when 493 => instruction_out <= x"00000003";
                when 494 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 495 => instruction_out <= x"040087c0";
                when 496 => instruction_out <= x"a0101003";   -- SSY 0x808;
                when 497 => instruction_out <= x"00000780";
                when 498 => instruction_out <= x"100fc003";   -- BRA (C48.EQU), 0x7e0;
                when 499 => instruction_out <= x"00000500";
                when 500 => instruction_out <= x"f0000001";   -- NOP;
                when 501 => instruction_out <= x"e0000000";
                when 502 => instruction_out <= x"10100003";   -- BRA 0x800;
                when 503 => instruction_out <= x"00000780";
                when 504 => instruction_out <= x"f0000001";   -- NOP;
                when 505 => instruction_out <= x"e0000000";
                when 506 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 507 => instruction_out <= x"80c00780";
                when 508 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 509 => instruction_out <= x"00000003";
                when 510 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 511 => instruction_out <= x"a0c00780";
                when 512 => instruction_out <= x"f0000001";   -- NOP;
                when 513 => instruction_out <= x"e0000000";
                when 514 => instruction_out <= x"f0000001";   -- NOP.S;
                when 515 => instruction_out <= x"e0000002";
                when 516 => instruction_out <= x"1015802d";   -- MVI R11, 0x15;
                when 517 => instruction_out <= x"00000003";
                when 518 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 519 => instruction_out <= x"040087c0";
                when 520 => instruction_out <= x"a010d003";   -- SSY 0x868;
                when 521 => instruction_out <= x"00000780";
                when 522 => instruction_out <= x"10108003";   -- BRA (C48.EQU), 0x840;
                when 523 => instruction_out <= x"00000500";
                when 524 => instruction_out <= x"f0000001";   -- NOP;
                when 525 => instruction_out <= x"e0000000";
                when 526 => instruction_out <= x"1010c003";   -- BRA 0x860;
                when 527 => instruction_out <= x"00000780";
                when 528 => instruction_out <= x"f0000001";   -- NOP;
                when 529 => instruction_out <= x"e0000000";
                when 530 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 531 => instruction_out <= x"80c00780";
                when 532 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 533 => instruction_out <= x"00000003";
                when 534 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 535 => instruction_out <= x"a0c00780";
                when 536 => instruction_out <= x"f0000001";   -- NOP;
                when 537 => instruction_out <= x"e0000000";
                when 538 => instruction_out <= x"f0000001";   -- NOP.S;
                when 539 => instruction_out <= x"e0000002";
                when 540 => instruction_out <= x"1016802d";   -- MVI R11, 0x16;
                when 541 => instruction_out <= x"00000003";
                when 542 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 543 => instruction_out <= x"040087c0";
                when 544 => instruction_out <= x"a0119003";   -- SSY 0x8c8;
                when 545 => instruction_out <= x"00000780";
                when 546 => instruction_out <= x"10114003";   -- BRA (C48.EQU), 0x8a0;
                when 547 => instruction_out <= x"00000500";
                when 548 => instruction_out <= x"f0000001";   -- NOP;
                when 549 => instruction_out <= x"e0000000";
                when 550 => instruction_out <= x"10118003";   -- BRA 0x8c0;
                when 551 => instruction_out <= x"00000780";
                when 552 => instruction_out <= x"f0000001";   -- NOP;
                when 553 => instruction_out <= x"e0000000";
                when 554 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 555 => instruction_out <= x"80c00780";
                when 556 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 557 => instruction_out <= x"00000003";
                when 558 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 559 => instruction_out <= x"a0c00780";
                when 560 => instruction_out <= x"f0000001";   -- NOP;
                when 561 => instruction_out <= x"e0000000";
                when 562 => instruction_out <= x"f0000001";   -- NOP.S;
                when 563 => instruction_out <= x"e0000002";
                when 564 => instruction_out <= x"1017802d";   -- MVI R11, 0x17;
                when 565 => instruction_out <= x"00000003";
                when 566 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 567 => instruction_out <= x"040087c0";
                when 568 => instruction_out <= x"a0125003";   -- SSY 0x928;
                when 569 => instruction_out <= x"00000780";
                when 570 => instruction_out <= x"10120003";   -- BRA (C48.EQU), 0x900;
                when 571 => instruction_out <= x"00000500";
                when 572 => instruction_out <= x"f0000001";   -- NOP;
                when 573 => instruction_out <= x"e0000000";
                when 574 => instruction_out <= x"10124003";   -- BRA 0x920;
                when 575 => instruction_out <= x"00000780";
                when 576 => instruction_out <= x"f0000001";   -- NOP;
                when 577 => instruction_out <= x"e0000000";
                when 578 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 579 => instruction_out <= x"80c00780";
                when 580 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 581 => instruction_out <= x"00000003";
                when 582 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 583 => instruction_out <= x"a0c00780";
                when 584 => instruction_out <= x"f0000001";   -- NOP;
                when 585 => instruction_out <= x"e0000000";
                when 586 => instruction_out <= x"f0000001";   -- NOP.S;
                when 587 => instruction_out <= x"e0000002";
                when 588 => instruction_out <= x"1018802d";   -- MVI R11, 0x18;
                when 589 => instruction_out <= x"00000003";
                when 590 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 591 => instruction_out <= x"040087c0";
                when 592 => instruction_out <= x"a0131003";   -- SSY 0x988;
                when 593 => instruction_out <= x"00000780";
                when 594 => instruction_out <= x"1012c003";   -- BRA (C48.EQU), 0x960;
                when 595 => instruction_out <= x"00000500";
                when 596 => instruction_out <= x"f0000001";   -- NOP;
                when 597 => instruction_out <= x"e0000000";
                when 598 => instruction_out <= x"10130003";   -- BRA 0x980;
                when 599 => instruction_out <= x"00000780";
                when 600 => instruction_out <= x"f0000001";   -- NOP;
                when 601 => instruction_out <= x"e0000000";
                when 602 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 603 => instruction_out <= x"80c00780";
                when 604 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 605 => instruction_out <= x"00000003";
                when 606 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 607 => instruction_out <= x"a0c00780";
                when 608 => instruction_out <= x"f0000001";   -- NOP;
                when 609 => instruction_out <= x"e0000000";
                when 610 => instruction_out <= x"f0000001";   -- NOP.S;
                when 611 => instruction_out <= x"e0000002";
                when 612 => instruction_out <= x"1019802d";   -- MVI R11, 0x19;
                when 613 => instruction_out <= x"00000003";
                when 614 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 615 => instruction_out <= x"040087c0";
                when 616 => instruction_out <= x"a013d003";   -- SSY 0x9e8;
                when 617 => instruction_out <= x"00000780";
                when 618 => instruction_out <= x"10138003";   -- BRA (C48.EQU), 0x9c0;
                when 619 => instruction_out <= x"00000500";
                when 620 => instruction_out <= x"f0000001";   -- NOP;
                when 621 => instruction_out <= x"e0000000";
                when 622 => instruction_out <= x"1013c003";   -- BRA 0x9e0;
                when 623 => instruction_out <= x"00000780";
                when 624 => instruction_out <= x"f0000001";   -- NOP;
                when 625 => instruction_out <= x"e0000000";
                when 626 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 627 => instruction_out <= x"80c00780";
                when 628 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 629 => instruction_out <= x"00000003";
                when 630 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 631 => instruction_out <= x"a0c00780";
                when 632 => instruction_out <= x"f0000001";   -- NOP;
                when 633 => instruction_out <= x"e0000000";
                when 634 => instruction_out <= x"f0000001";   -- NOP.S;
                when 635 => instruction_out <= x"e0000002";
                when 636 => instruction_out <= x"101a802d";   -- MVI R11, 0x1a;
                when 637 => instruction_out <= x"00000003";
                when 638 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 639 => instruction_out <= x"040087c0";
                when 640 => instruction_out <= x"a0149003";   -- SSY 0xa48;
                when 641 => instruction_out <= x"00000780";
                when 642 => instruction_out <= x"10144003";   -- BRA (C48.EQU), 0xa20;
                when 643 => instruction_out <= x"00000500";
                when 644 => instruction_out <= x"f0000001";   -- NOP;
                when 645 => instruction_out <= x"e0000000";
                when 646 => instruction_out <= x"10148003";   -- BRA 0xa40;
                when 647 => instruction_out <= x"00000780";
                when 648 => instruction_out <= x"f0000001";   -- NOP;
                when 649 => instruction_out <= x"e0000000";
                when 650 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 651 => instruction_out <= x"80c00780";
                when 652 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 653 => instruction_out <= x"00000003";
                when 654 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 655 => instruction_out <= x"a0c00780";
                when 656 => instruction_out <= x"f0000001";   -- NOP;
                when 657 => instruction_out <= x"e0000000";
                when 658 => instruction_out <= x"f0000001";   -- NOP.S;
                when 659 => instruction_out <= x"e0000002";
                when 660 => instruction_out <= x"101b802d";   -- MVI R11, 0x1b;
                when 661 => instruction_out <= x"00000003";
                when 662 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 663 => instruction_out <= x"040087c0";
                when 664 => instruction_out <= x"a0155003";   -- SSY 0xaa8;
                when 665 => instruction_out <= x"00000780";
                when 666 => instruction_out <= x"10150003";   -- BRA (C48.EQU), 0xa80;
                when 667 => instruction_out <= x"00000500";
                when 668 => instruction_out <= x"f0000001";   -- NOP;
                when 669 => instruction_out <= x"e0000000";
                when 670 => instruction_out <= x"10154003";   -- BRA 0xaa0;
                when 671 => instruction_out <= x"00000780";
                when 672 => instruction_out <= x"f0000001";   -- NOP;
                when 673 => instruction_out <= x"e0000000";
                when 674 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 675 => instruction_out <= x"80c00780";
                when 676 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 677 => instruction_out <= x"00000003";
                when 678 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 679 => instruction_out <= x"a0c00780";
                when 680 => instruction_out <= x"f0000001";   -- NOP;
                when 681 => instruction_out <= x"e0000000";
                when 682 => instruction_out <= x"f0000001";   -- NOP.S;
                when 683 => instruction_out <= x"e0000002";
                when 684 => instruction_out <= x"101c802d";   -- MVI R11, 0x1c;
                when 685 => instruction_out <= x"00000003";
                when 686 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 687 => instruction_out <= x"040087c0";
                when 688 => instruction_out <= x"a0161003";   -- SSY 0xb08;
                when 689 => instruction_out <= x"00000780";
                when 690 => instruction_out <= x"1015c003";   -- BRA (C48.EQU), 0xae0;
                when 691 => instruction_out <= x"00000500";
                when 692 => instruction_out <= x"f0000001";   -- NOP;
                when 693 => instruction_out <= x"e0000000";
                when 694 => instruction_out <= x"10160003";   -- BRA 0xb00;
                when 695 => instruction_out <= x"00000780";
                when 696 => instruction_out <= x"f0000001";   -- NOP;
                when 697 => instruction_out <= x"e0000000";
                when 698 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 699 => instruction_out <= x"80c00780";
                when 700 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 701 => instruction_out <= x"00000003";
                when 702 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 703 => instruction_out <= x"a0c00780";
                when 704 => instruction_out <= x"f0000001";   -- NOP;
                when 705 => instruction_out <= x"e0000000";
                when 706 => instruction_out <= x"f0000001";   -- NOP.S;
                when 707 => instruction_out <= x"e0000002";
                when 708 => instruction_out <= x"101d802d";   -- MVI R11, 0x1d;
                when 709 => instruction_out <= x"00000003";
                when 710 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 711 => instruction_out <= x"040087c0";
                when 712 => instruction_out <= x"a016d003";   -- SSY 0xb68;
                when 713 => instruction_out <= x"00000780";
                when 714 => instruction_out <= x"10168003";   -- BRA (C48.EQU), 0xb40;
                when 715 => instruction_out <= x"00000500";
                when 716 => instruction_out <= x"f0000001";   -- NOP;
                when 717 => instruction_out <= x"e0000000";
                when 718 => instruction_out <= x"1016c003";   -- BRA 0xb60;
                when 719 => instruction_out <= x"00000780";
                when 720 => instruction_out <= x"f0000001";   -- NOP;
                when 721 => instruction_out <= x"e0000000";
                when 722 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 723 => instruction_out <= x"80c00780";
                when 724 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 725 => instruction_out <= x"00000003";
                when 726 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 727 => instruction_out <= x"a0c00780";
                when 728 => instruction_out <= x"f0000001";   -- NOP;
                when 729 => instruction_out <= x"e0000000";
                when 730 => instruction_out <= x"f0000001";   -- NOP.S;
                when 731 => instruction_out <= x"e0000002";
                when 732 => instruction_out <= x"101e802d";   -- MVI R11, 0x1e;
                when 733 => instruction_out <= x"00000003";
                when 734 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 735 => instruction_out <= x"040087c0";
                when 736 => instruction_out <= x"a0179003";   -- SSY 0xbc8;
                when 737 => instruction_out <= x"00000780";
                when 738 => instruction_out <= x"10174003";   -- BRA (C48.EQU), 0xba0;
                when 739 => instruction_out <= x"00000500";
                when 740 => instruction_out <= x"f0000001";   -- NOP;
                when 741 => instruction_out <= x"e0000000";
                when 742 => instruction_out <= x"10178003";   -- BRA 0xbc0;
                when 743 => instruction_out <= x"00000780";
                when 744 => instruction_out <= x"f0000001";   -- NOP;
                when 745 => instruction_out <= x"e0000000";
                when 746 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 747 => instruction_out <= x"80c00780";
                when 748 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 749 => instruction_out <= x"00000003";
                when 750 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 751 => instruction_out <= x"a0c00780";
                when 752 => instruction_out <= x"f0000001";   -- NOP;
                when 753 => instruction_out <= x"e0000000";
                when 754 => instruction_out <= x"f0000001";   -- NOP.S;
                when 755 => instruction_out <= x"e0000002";
                when 756 => instruction_out <= x"101f802d";   -- MVI R11, 0x1f;
                when 757 => instruction_out <= x"00000003";
                when 758 => instruction_out <= x"d00a1639";   -- LOP.XOR.C0 R14, R11, R10;
                when 759 => instruction_out <= x"040087c0";
                when 760 => instruction_out <= x"a0185003";   -- SSY 0xc28;
                when 761 => instruction_out <= x"00000780";
                when 762 => instruction_out <= x"10180003";   -- BRA (C48.EQU), 0xc00;
                when 763 => instruction_out <= x"00000500";
                when 764 => instruction_out <= x"f0000001";   -- NOP;
                when 765 => instruction_out <= x"e0000000";
                when 766 => instruction_out <= x"10184003";   -- BRA 0xc20;
                when 767 => instruction_out <= x"00000780";
                when 768 => instruction_out <= x"f0000001";   -- NOP;
                when 769 => instruction_out <= x"e0000000";
                when 770 => instruction_out <= x"d00e1835";   -- GLD.U32 R13, global14 [R12];
                when 771 => instruction_out <= x"80c00780";
                when 772 => instruction_out <= x"20019a35";   -- IADD32I R13, R13, 0x1;
                when 773 => instruction_out <= x"00000003";
                when 774 => instruction_out <= x"d00e1835";   -- GST.U32 global14 [R12], R13;
                when 775 => instruction_out <= x"a0c00780";
                when 776 => instruction_out <= x"f0000001";   -- NOP;
                when 777 => instruction_out <= x"e0000000";
                when 778 => instruction_out <= x"f0000001";   -- NOP.S;
                when 779 => instruction_out <= x"e0000002";
                when 780 => instruction_out <= x"30000003";   -- RET;
                when 781 => instruction_out <= x"00000780";
                when 782 => instruction_out <= x"f0000001";   -- NOP;
                when 783 => instruction_out <= x"e0000000";
                when 784 => instruction_out <= x"30000003";   -- RET
                when 785 => instruction_out <= x"00000780";

			when others => null;
		end case;
	end process;

end arch;

